////////////////////////////////////////////////////////////////////////////
// Author       : Prajyot 
// Coursework   : ECE 751
// Module       : adder_tree
// Description  : Adder tree logic, which takes in the tlut prodict matrix
//                and add relevant indexes to provide the matrix
//                multiplication results. Generated using gen.cpp file
////////////////////////////////////////////////////////////////////////////

`include "DEF.sv"
module adder_tree(
    input  logic clk,
    input  logic rst_n,
    input  logic [`DIM_ROW2 * `DIM_COL2 -1:0][`DIM_ROW1 * `DIM_COL1 -1:0][`ACC_WIDTH-1:0]prod,
    output logic [`DIM_ROW1 * `DIM_COL2 -1:0][`ACC_WIDTH-1:0]mult
    //TODO: Update the DIM of the output
    //for now, it is = DIM_A
    //Aish: Changed DIM_A = DIM_ROW1 * DIM_COL1
    //Aish: Changed DIM_C = DIM_ROW2 * DIM_COL2
    //Aish: Changed DIM_MULT = DIM_ROW1 * DIM_COL2
);
    logic [`DIM_ROW1 * `DIM_COL2 -1:0][`ACC_WIDTH-1:0] mul_temp;

    always_ff @(posedge clk or negedge rst_n)
    begin
        if(~rst_n)
            mul_temp <= 0;
        else
        begin
        // Below code generated using ./_gen_add_logic <array dim> 
mul_temp[0] = prod[0][0] + prod[1][10] + prod[2][20] + prod[3][30] + prod[4][40] + prod[5][50] + prod[6][60] + prod[7][70] + prod[8][80] + prod[9][90] + prod[10][100] + prod[11][110] + prod[12][120] + prod[13][130] + prod[14][140] + prod[15][150] + prod[16][160] + prod[17][170] + prod[18][180] + prod[19][190] + prod[20][200] + prod[21][210] + prod[22][220] + prod[23][230] + prod[24][240] + prod[25][250] + prod[26][260] + prod[27][270] + prod[28][280] + prod[29][290] + prod[30][300] + prod[31][310] + prod[32][320] + prod[33][330] + prod[34][340] + prod[35][350] + prod[36][360] + prod[37][370] + prod[38][380] + prod[39][390] + prod[40][400] + prod[41][410] + prod[42][420] + prod[43][430] + prod[44][440] + prod[45][450] + prod[46][460] + prod[47][470] + prod[48][480] + prod[49][490] + prod[50][500] + prod[51][510] + prod[52][520] + prod[53][530] + prod[54][540] + prod[55][550] + prod[56][560] + prod[57][570] + prod[58][580] + prod[59][590] + prod[60][600] + prod[61][610] + prod[62][620] + prod[63][630] + prod[64][640] + prod[65][650] + prod[66][660] + prod[67][670] + prod[68][680] + prod[69][690] + prod[70][700] + prod[71][710] + prod[72][720] + prod[73][730] + prod[74][740] + prod[75][750] + prod[76][760] + prod[77][770] + prod[78][780] + prod[79][790] + prod[80][800] + prod[81][810] + prod[82][820] + prod[83][830] + prod[84][840] + prod[85][850] + prod[86][860] + prod[87][870] + prod[88][880] + prod[89][890] + prod[90][900] + prod[91][910] + prod[92][920] + prod[93][930] + prod[94][940] + prod[95][950] + prod[96][960] + prod[97][970] + prod[98][980] + prod[99][990] + prod[100][1000] + prod[101][1010] + prod[102][1020] + prod[103][1030] + prod[104][1040] + prod[105][1050] + prod[106][1060] + prod[107][1070] + prod[108][1080] + prod[109][1090] + prod[110][1100] + prod[111][1110] + prod[112][1120] + prod[113][1130] + prod[114][1140] + prod[115][1150] + prod[116][1160] + prod[117][1170] + prod[118][1180] + prod[119][1190] + prod[120][1200] + prod[121][1210] + prod[122][1220] + prod[123][1230] + prod[124][1240] + prod[125][1250] + prod[126][1260] + prod[127][1270] + prod[128][1280] + prod[129][1290] + prod[130][1300] + prod[131][1310] + prod[132][1320] + prod[133][1330] + prod[134][1340] + prod[135][1350] + prod[136][1360] + prod[137][1370] + prod[138][1380] + prod[139][1390] + prod[140][1400] + prod[141][1410] + prod[142][1420] + prod[143][1430] + prod[144][1440] + prod[145][1450] + prod[146][1460] + prod[147][1470] + prod[148][1480] + prod[149][1490] + prod[150][1500] + prod[151][1510] + prod[152][1520] + prod[153][1530] + prod[154][1540] + prod[155][1550] + prod[156][1560] + prod[157][1570] + prod[158][1580] + prod[159][1590] + prod[160][1600] + prod[161][1610] + prod[162][1620] + prod[163][1630] + prod[164][1640] + prod[165][1650] + prod[166][1660] + prod[167][1670] + prod[168][1680] + prod[169][1690] + prod[170][1700] + prod[171][1710] + prod[172][1720] + prod[173][1730] + prod[174][1740] + prod[175][1750] + prod[176][1760] + prod[177][1770] + prod[178][1780] + prod[179][1790] + prod[180][1800] + prod[181][1810] + prod[182][1820] + prod[183][1830] + prod[184][1840] + prod[185][1850] + prod[186][1860] + prod[187][1870] + prod[188][1880] + prod[189][1890] + prod[190][1900] + prod[191][1910] + prod[192][1920] + prod[193][1930] + prod[194][1940] + prod[195][1950] + prod[196][1960] + prod[197][1970] + prod[198][1980] + prod[199][1990] + prod[200][2000] + prod[201][2010] + prod[202][2020] + prod[203][2030] + prod[204][2040] + prod[205][2050] + prod[206][2060] + prod[207][2070] + prod[208][2080] + prod[209][2090] + prod[210][2100] + prod[211][2110] + prod[212][2120] + prod[213][2130] + prod[214][2140] + prod[215][2150] + prod[216][2160] + prod[217][2170] + prod[218][2180] + prod[219][2190] + prod[220][2200] + prod[221][2210] + prod[222][2220] + prod[223][2230] + prod[224][2240] + prod[225][2250] + prod[226][2260] + prod[227][2270] + prod[228][2280] + prod[229][2290] + prod[230][2300] + prod[231][2310] + prod[232][2320] + prod[233][2330] + prod[234][2340] + prod[235][2350] + prod[236][2360] + prod[237][2370] + prod[238][2380] + prod[239][2390] + prod[240][2400] + prod[241][2410] + prod[242][2420] + prod[243][2430] + prod[244][2440] + prod[245][2450] + prod[246][2460] + prod[247][2470] + prod[248][2480] + prod[249][2490] + prod[250][2500] + prod[251][2510] + prod[252][2520] + prod[253][2530] + prod[254][2540] + prod[255][2550] + prod[256][2560] + prod[257][2570] + prod[258][2580] + prod[259][2590] + prod[260][2600] + prod[261][2610] + prod[262][2620] + prod[263][2630] + prod[264][2640] + prod[265][2650] + prod[266][2660] + prod[267][2670] + prod[268][2680] + prod[269][2690] + prod[270][2700] + prod[271][2710] + prod[272][2720] + prod[273][2730] + prod[274][2740] + prod[275][2750] + prod[276][2760] + prod[277][2770] + prod[278][2780] + prod[279][2790] + prod[280][2800] + prod[281][2810] + prod[282][2820] + prod[283][2830] + prod[284][2840] + prod[285][2850] + prod[286][2860] + prod[287][2870] + prod[288][2880] + prod[289][2890] + prod[290][2900] + prod[291][2910] + prod[292][2920] + prod[293][2930] + prod[294][2940] + prod[295][2950] + prod[296][2960] + prod[297][2970] + prod[298][2980] + prod[299][2990] + prod[300][3000] + prod[301][3010] + prod[302][3020] + prod[303][3030] + prod[304][3040] + prod[305][3050] + prod[306][3060] + prod[307][3070] + prod[308][3080] + prod[309][3090] + prod[310][3100] + prod[311][3110] + prod[312][3120] + prod[313][3130] + prod[314][3140] + prod[315][3150] + prod[316][3160] + prod[317][3170] + prod[318][3180] + prod[319][3190] + prod[320][3200] + prod[321][3210] + prod[322][3220] + prod[323][3230] + prod[324][3240] + prod[325][3250] + prod[326][3260] + prod[327][3270] + prod[328][3280] + prod[329][3290] + prod[330][3300] + prod[331][3310] + prod[332][3320] + prod[333][3330] + prod[334][3340] + prod[335][3350] + prod[336][3360] + prod[337][3370] + prod[338][3380] + prod[339][3390] + prod[340][3400] + prod[341][3410] + prod[342][3420] + prod[343][3430] + prod[344][3440] + prod[345][3450] + prod[346][3460] + prod[347][3470] + prod[348][3480] + prod[349][3490] + prod[350][3500] + prod[351][3510] + prod[352][3520] + prod[353][3530] + prod[354][3540] + prod[355][3550] + prod[356][3560] + prod[357][3570] + prod[358][3580] + prod[359][3590] + prod[360][3600] + prod[361][3610] + prod[362][3620] + prod[363][3630] + prod[364][3640] + prod[365][3650] + prod[366][3660] + prod[367][3670] + prod[368][3680] + prod[369][3690] + prod[370][3700] + prod[371][3710] + prod[372][3720] + prod[373][3730] + prod[374][3740] + prod[375][3750] + prod[376][3760] + prod[377][3770] + prod[378][3780] + prod[379][3790] + prod[380][3800] + prod[381][3810] + prod[382][3820] + prod[383][3830] + prod[384][3840] + prod[385][3850] + prod[386][3860] + prod[387][3870] + prod[388][3880] + prod[389][3890] + prod[390][3900] + prod[391][3910] + prod[392][3920] + prod[393][3930] + prod[394][3940] + prod[395][3950] + prod[396][3960] + prod[397][3970] + prod[398][3980] + prod[399][3990] + prod[400][4000] + prod[401][4010] + prod[402][4020] + prod[403][4030] + prod[404][4040] + prod[405][4050] + prod[406][4060] + prod[407][4070] + prod[408][4080] + prod[409][4090] + prod[410][4100] + prod[411][4110] + prod[412][4120] + prod[413][4130] + prod[414][4140] + prod[415][4150] + prod[416][4160] + prod[417][4170] + prod[418][4180] + prod[419][4190] + prod[420][4200] + prod[421][4210] + prod[422][4220] + prod[423][4230] + prod[424][4240] + prod[425][4250] + prod[426][4260] + prod[427][4270] + prod[428][4280] + prod[429][4290] + prod[430][4300] + prod[431][4310] + prod[432][4320] + prod[433][4330] + prod[434][4340] + prod[435][4350] + prod[436][4360] + prod[437][4370] + prod[438][4380] + prod[439][4390] + prod[440][4400] + prod[441][4410] + prod[442][4420] + prod[443][4430] + prod[444][4440] + prod[445][4450] + prod[446][4460] + prod[447][4470] + prod[448][4480] + prod[449][4490] + prod[450][4500] + prod[451][4510] + prod[452][4520] + prod[453][4530] + prod[454][4540] + prod[455][4550] + prod[456][4560] + prod[457][4570] + prod[458][4580] + prod[459][4590] + prod[460][4600] + prod[461][4610] + prod[462][4620] + prod[463][4630] + prod[464][4640] + prod[465][4650] + prod[466][4660] + prod[467][4670] + prod[468][4680] + prod[469][4690] + prod[470][4700] + prod[471][4710] + prod[472][4720] + prod[473][4730] + prod[474][4740] + prod[475][4750] + prod[476][4760] + prod[477][4770] + prod[478][4780] + prod[479][4790] + prod[480][4800] + prod[481][4810] + prod[482][4820] + prod[483][4830] + prod[484][4840] + prod[485][4850] + prod[486][4860] + prod[487][4870] + prod[488][4880] + prod[489][4890] + prod[490][4900] + prod[491][4910] + prod[492][4920] + prod[493][4930] + prod[494][4940] + prod[495][4950] + prod[496][4960] + prod[497][4970] + prod[498][4980] + prod[499][4990] + prod[500][5000] + prod[501][5010] + prod[502][5020] + prod[503][5030] + prod[504][5040] + prod[505][5050] + prod[506][5060] + prod[507][5070] + prod[508][5080] + prod[509][5090] + prod[510][5100] + prod[511][5110] + prod[512][5120] + prod[513][5130] + prod[514][5140] + prod[515][5150] + prod[516][5160] + prod[517][5170] + prod[518][5180] + prod[519][5190] + prod[520][5200] + prod[521][5210] + prod[522][5220] + prod[523][5230] + prod[524][5240] + prod[525][5250] + prod[526][5260] + prod[527][5270] + prod[528][5280] + prod[529][5290] + prod[530][5300] + prod[531][5310] + prod[532][5320] + prod[533][5330] + prod[534][5340] + prod[535][5350] + prod[536][5360] + prod[537][5370] + prod[538][5380] + prod[539][5390] + prod[540][5400] + prod[541][5410] + prod[542][5420] + prod[543][5430] + prod[544][5440] + prod[545][5450] + prod[546][5460] + prod[547][5470] + prod[548][5480] + prod[549][5490] + prod[550][5500] + prod[551][5510] + prod[552][5520] + prod[553][5530] + prod[554][5540] + prod[555][5550] + prod[556][5560] + prod[557][5570] + prod[558][5580] + prod[559][5590] + prod[560][5600] + prod[561][5610] + prod[562][5620] + prod[563][5630] + prod[564][5640] + prod[565][5650] + prod[566][5660] + prod[567][5670] + prod[568][5680] + prod[569][5690] + prod[570][5700] + prod[571][5710] + prod[572][5720] + prod[573][5730] + prod[574][5740] + prod[575][5750] + prod[576][5760] + prod[577][5770] + prod[578][5780] + prod[579][5790] + prod[580][5800] + prod[581][5810] + prod[582][5820] + prod[583][5830] + prod[584][5840] + prod[585][5850] + prod[586][5860] + prod[587][5870] + prod[588][5880] + prod[589][5890] + prod[590][5900] + prod[591][5910] + prod[592][5920] + prod[593][5930] + prod[594][5940] + prod[595][5950] + prod[596][5960] + prod[597][5970] + prod[598][5980] + prod[599][5990] + prod[600][6000] + prod[601][6010] + prod[602][6020] + prod[603][6030] + prod[604][6040] + prod[605][6050] + prod[606][6060] + prod[607][6070] + prod[608][6080] + prod[609][6090] + prod[610][6100] + prod[611][6110] + prod[612][6120] + prod[613][6130] + prod[614][6140] + prod[615][6150] + prod[616][6160] + prod[617][6170] + prod[618][6180] + prod[619][6190] + prod[620][6200] + prod[621][6210] + prod[622][6220] + prod[623][6230] + prod[624][6240] + prod[625][6250] + prod[626][6260] + prod[627][6270] + prod[628][6280] + prod[629][6290] + prod[630][6300] + prod[631][6310] + prod[632][6320] + prod[633][6330] + prod[634][6340] + prod[635][6350] + prod[636][6360] + prod[637][6370] + prod[638][6380] + prod[639][6390] + prod[640][6400] + prod[641][6410] + prod[642][6420] + prod[643][6430] + prod[644][6440] + prod[645][6450] + prod[646][6460] + prod[647][6470] + prod[648][6480] + prod[649][6490] + prod[650][6500] + prod[651][6510] + prod[652][6520] + prod[653][6530] + prod[654][6540] + prod[655][6550] + prod[656][6560] + prod[657][6570] + prod[658][6580] + prod[659][6590] + prod[660][6600] + prod[661][6610] + prod[662][6620] + prod[663][6630] + prod[664][6640] + prod[665][6650] + prod[666][6660] + prod[667][6670] + prod[668][6680] + prod[669][6690] + prod[670][6700] + prod[671][6710] + prod[672][6720] + prod[673][6730] + prod[674][6740] + prod[675][6750] + prod[676][6760] + prod[677][6770] + prod[678][6780] + prod[679][6790] + prod[680][6800] + prod[681][6810] + prod[682][6820] + prod[683][6830] + prod[684][6840] + prod[685][6850] + prod[686][6860] + prod[687][6870] + prod[688][6880] + prod[689][6890] + prod[690][6900] + prod[691][6910] + prod[692][6920] + prod[693][6930] + prod[694][6940] + prod[695][6950] + prod[696][6960] + prod[697][6970] + prod[698][6980] + prod[699][6990] + prod[700][7000] + prod[701][7010] + prod[702][7020] + prod[703][7030] + prod[704][7040] + prod[705][7050] + prod[706][7060] + prod[707][7070] + prod[708][7080] + prod[709][7090] + prod[710][7100] + prod[711][7110] + prod[712][7120] + prod[713][7130] + prod[714][7140] + prod[715][7150] + prod[716][7160] + prod[717][7170] + prod[718][7180] + prod[719][7190] + prod[720][7200] + prod[721][7210] + prod[722][7220] + prod[723][7230] + prod[724][7240] + prod[725][7250] + prod[726][7260] + prod[727][7270] + prod[728][7280] + prod[729][7290] + prod[730][7300] + prod[731][7310] + prod[732][7320] + prod[733][7330] + prod[734][7340] + prod[735][7350] + prod[736][7360] + prod[737][7370] + prod[738][7380] + prod[739][7390] + prod[740][7400] + prod[741][7410] + prod[742][7420] + prod[743][7430] + prod[744][7440] + prod[745][7450] + prod[746][7460] + prod[747][7470] + prod[748][7480] + prod[749][7490] + prod[750][7500] + prod[751][7510] + prod[752][7520] + prod[753][7530] + prod[754][7540] + prod[755][7550] + prod[756][7560] + prod[757][7570] + prod[758][7580] + prod[759][7590] + prod[760][7600] + prod[761][7610] + prod[762][7620] + prod[763][7630] + prod[764][7640] + prod[765][7650] + prod[766][7660] + prod[767][7670] + prod[768][7680] + prod[769][7690] + prod[770][7700] + prod[771][7710] + prod[772][7720] + prod[773][7730] + prod[774][7740] + prod[775][7750] + prod[776][7760] + prod[777][7770] + prod[778][7780] + prod[779][7790] + prod[780][7800] + prod[781][7810] + prod[782][7820] + prod[783][7830];
mul_temp[1] = prod[0][1] + prod[1][11] + prod[2][21] + prod[3][31] + prod[4][41] + prod[5][51] + prod[6][61] + prod[7][71] + prod[8][81] + prod[9][91] + prod[10][101] + prod[11][111] + prod[12][121] + prod[13][131] + prod[14][141] + prod[15][151] + prod[16][161] + prod[17][171] + prod[18][181] + prod[19][191] + prod[20][201] + prod[21][211] + prod[22][221] + prod[23][231] + prod[24][241] + prod[25][251] + prod[26][261] + prod[27][271] + prod[28][281] + prod[29][291] + prod[30][301] + prod[31][311] + prod[32][321] + prod[33][331] + prod[34][341] + prod[35][351] + prod[36][361] + prod[37][371] + prod[38][381] + prod[39][391] + prod[40][401] + prod[41][411] + prod[42][421] + prod[43][431] + prod[44][441] + prod[45][451] + prod[46][461] + prod[47][471] + prod[48][481] + prod[49][491] + prod[50][501] + prod[51][511] + prod[52][521] + prod[53][531] + prod[54][541] + prod[55][551] + prod[56][561] + prod[57][571] + prod[58][581] + prod[59][591] + prod[60][601] + prod[61][611] + prod[62][621] + prod[63][631] + prod[64][641] + prod[65][651] + prod[66][661] + prod[67][671] + prod[68][681] + prod[69][691] + prod[70][701] + prod[71][711] + prod[72][721] + prod[73][731] + prod[74][741] + prod[75][751] + prod[76][761] + prod[77][771] + prod[78][781] + prod[79][791] + prod[80][801] + prod[81][811] + prod[82][821] + prod[83][831] + prod[84][841] + prod[85][851] + prod[86][861] + prod[87][871] + prod[88][881] + prod[89][891] + prod[90][901] + prod[91][911] + prod[92][921] + prod[93][931] + prod[94][941] + prod[95][951] + prod[96][961] + prod[97][971] + prod[98][981] + prod[99][991] + prod[100][1001] + prod[101][1011] + prod[102][1021] + prod[103][1031] + prod[104][1041] + prod[105][1051] + prod[106][1061] + prod[107][1071] + prod[108][1081] + prod[109][1091] + prod[110][1101] + prod[111][1111] + prod[112][1121] + prod[113][1131] + prod[114][1141] + prod[115][1151] + prod[116][1161] + prod[117][1171] + prod[118][1181] + prod[119][1191] + prod[120][1201] + prod[121][1211] + prod[122][1221] + prod[123][1231] + prod[124][1241] + prod[125][1251] + prod[126][1261] + prod[127][1271] + prod[128][1281] + prod[129][1291] + prod[130][1301] + prod[131][1311] + prod[132][1321] + prod[133][1331] + prod[134][1341] + prod[135][1351] + prod[136][1361] + prod[137][1371] + prod[138][1381] + prod[139][1391] + prod[140][1401] + prod[141][1411] + prod[142][1421] + prod[143][1431] + prod[144][1441] + prod[145][1451] + prod[146][1461] + prod[147][1471] + prod[148][1481] + prod[149][1491] + prod[150][1501] + prod[151][1511] + prod[152][1521] + prod[153][1531] + prod[154][1541] + prod[155][1551] + prod[156][1561] + prod[157][1571] + prod[158][1581] + prod[159][1591] + prod[160][1601] + prod[161][1611] + prod[162][1621] + prod[163][1631] + prod[164][1641] + prod[165][1651] + prod[166][1661] + prod[167][1671] + prod[168][1681] + prod[169][1691] + prod[170][1701] + prod[171][1711] + prod[172][1721] + prod[173][1731] + prod[174][1741] + prod[175][1751] + prod[176][1761] + prod[177][1771] + prod[178][1781] + prod[179][1791] + prod[180][1801] + prod[181][1811] + prod[182][1821] + prod[183][1831] + prod[184][1841] + prod[185][1851] + prod[186][1861] + prod[187][1871] + prod[188][1881] + prod[189][1891] + prod[190][1901] + prod[191][1911] + prod[192][1921] + prod[193][1931] + prod[194][1941] + prod[195][1951] + prod[196][1961] + prod[197][1971] + prod[198][1981] + prod[199][1991] + prod[200][2001] + prod[201][2011] + prod[202][2021] + prod[203][2031] + prod[204][2041] + prod[205][2051] + prod[206][2061] + prod[207][2071] + prod[208][2081] + prod[209][2091] + prod[210][2101] + prod[211][2111] + prod[212][2121] + prod[213][2131] + prod[214][2141] + prod[215][2151] + prod[216][2161] + prod[217][2171] + prod[218][2181] + prod[219][2191] + prod[220][2201] + prod[221][2211] + prod[222][2221] + prod[223][2231] + prod[224][2241] + prod[225][2251] + prod[226][2261] + prod[227][2271] + prod[228][2281] + prod[229][2291] + prod[230][2301] + prod[231][2311] + prod[232][2321] + prod[233][2331] + prod[234][2341] + prod[235][2351] + prod[236][2361] + prod[237][2371] + prod[238][2381] + prod[239][2391] + prod[240][2401] + prod[241][2411] + prod[242][2421] + prod[243][2431] + prod[244][2441] + prod[245][2451] + prod[246][2461] + prod[247][2471] + prod[248][2481] + prod[249][2491] + prod[250][2501] + prod[251][2511] + prod[252][2521] + prod[253][2531] + prod[254][2541] + prod[255][2551] + prod[256][2561] + prod[257][2571] + prod[258][2581] + prod[259][2591] + prod[260][2601] + prod[261][2611] + prod[262][2621] + prod[263][2631] + prod[264][2641] + prod[265][2651] + prod[266][2661] + prod[267][2671] + prod[268][2681] + prod[269][2691] + prod[270][2701] + prod[271][2711] + prod[272][2721] + prod[273][2731] + prod[274][2741] + prod[275][2751] + prod[276][2761] + prod[277][2771] + prod[278][2781] + prod[279][2791] + prod[280][2801] + prod[281][2811] + prod[282][2821] + prod[283][2831] + prod[284][2841] + prod[285][2851] + prod[286][2861] + prod[287][2871] + prod[288][2881] + prod[289][2891] + prod[290][2901] + prod[291][2911] + prod[292][2921] + prod[293][2931] + prod[294][2941] + prod[295][2951] + prod[296][2961] + prod[297][2971] + prod[298][2981] + prod[299][2991] + prod[300][3001] + prod[301][3011] + prod[302][3021] + prod[303][3031] + prod[304][3041] + prod[305][3051] + prod[306][3061] + prod[307][3071] + prod[308][3081] + prod[309][3091] + prod[310][3101] + prod[311][3111] + prod[312][3121] + prod[313][3131] + prod[314][3141] + prod[315][3151] + prod[316][3161] + prod[317][3171] + prod[318][3181] + prod[319][3191] + prod[320][3201] + prod[321][3211] + prod[322][3221] + prod[323][3231] + prod[324][3241] + prod[325][3251] + prod[326][3261] + prod[327][3271] + prod[328][3281] + prod[329][3291] + prod[330][3301] + prod[331][3311] + prod[332][3321] + prod[333][3331] + prod[334][3341] + prod[335][3351] + prod[336][3361] + prod[337][3371] + prod[338][3381] + prod[339][3391] + prod[340][3401] + prod[341][3411] + prod[342][3421] + prod[343][3431] + prod[344][3441] + prod[345][3451] + prod[346][3461] + prod[347][3471] + prod[348][3481] + prod[349][3491] + prod[350][3501] + prod[351][3511] + prod[352][3521] + prod[353][3531] + prod[354][3541] + prod[355][3551] + prod[356][3561] + prod[357][3571] + prod[358][3581] + prod[359][3591] + prod[360][3601] + prod[361][3611] + prod[362][3621] + prod[363][3631] + prod[364][3641] + prod[365][3651] + prod[366][3661] + prod[367][3671] + prod[368][3681] + prod[369][3691] + prod[370][3701] + prod[371][3711] + prod[372][3721] + prod[373][3731] + prod[374][3741] + prod[375][3751] + prod[376][3761] + prod[377][3771] + prod[378][3781] + prod[379][3791] + prod[380][3801] + prod[381][3811] + prod[382][3821] + prod[383][3831] + prod[384][3841] + prod[385][3851] + prod[386][3861] + prod[387][3871] + prod[388][3881] + prod[389][3891] + prod[390][3901] + prod[391][3911] + prod[392][3921] + prod[393][3931] + prod[394][3941] + prod[395][3951] + prod[396][3961] + prod[397][3971] + prod[398][3981] + prod[399][3991] + prod[400][4001] + prod[401][4011] + prod[402][4021] + prod[403][4031] + prod[404][4041] + prod[405][4051] + prod[406][4061] + prod[407][4071] + prod[408][4081] + prod[409][4091] + prod[410][4101] + prod[411][4111] + prod[412][4121] + prod[413][4131] + prod[414][4141] + prod[415][4151] + prod[416][4161] + prod[417][4171] + prod[418][4181] + prod[419][4191] + prod[420][4201] + prod[421][4211] + prod[422][4221] + prod[423][4231] + prod[424][4241] + prod[425][4251] + prod[426][4261] + prod[427][4271] + prod[428][4281] + prod[429][4291] + prod[430][4301] + prod[431][4311] + prod[432][4321] + prod[433][4331] + prod[434][4341] + prod[435][4351] + prod[436][4361] + prod[437][4371] + prod[438][4381] + prod[439][4391] + prod[440][4401] + prod[441][4411] + prod[442][4421] + prod[443][4431] + prod[444][4441] + prod[445][4451] + prod[446][4461] + prod[447][4471] + prod[448][4481] + prod[449][4491] + prod[450][4501] + prod[451][4511] + prod[452][4521] + prod[453][4531] + prod[454][4541] + prod[455][4551] + prod[456][4561] + prod[457][4571] + prod[458][4581] + prod[459][4591] + prod[460][4601] + prod[461][4611] + prod[462][4621] + prod[463][4631] + prod[464][4641] + prod[465][4651] + prod[466][4661] + prod[467][4671] + prod[468][4681] + prod[469][4691] + prod[470][4701] + prod[471][4711] + prod[472][4721] + prod[473][4731] + prod[474][4741] + prod[475][4751] + prod[476][4761] + prod[477][4771] + prod[478][4781] + prod[479][4791] + prod[480][4801] + prod[481][4811] + prod[482][4821] + prod[483][4831] + prod[484][4841] + prod[485][4851] + prod[486][4861] + prod[487][4871] + prod[488][4881] + prod[489][4891] + prod[490][4901] + prod[491][4911] + prod[492][4921] + prod[493][4931] + prod[494][4941] + prod[495][4951] + prod[496][4961] + prod[497][4971] + prod[498][4981] + prod[499][4991] + prod[500][5001] + prod[501][5011] + prod[502][5021] + prod[503][5031] + prod[504][5041] + prod[505][5051] + prod[506][5061] + prod[507][5071] + prod[508][5081] + prod[509][5091] + prod[510][5101] + prod[511][5111] + prod[512][5121] + prod[513][5131] + prod[514][5141] + prod[515][5151] + prod[516][5161] + prod[517][5171] + prod[518][5181] + prod[519][5191] + prod[520][5201] + prod[521][5211] + prod[522][5221] + prod[523][5231] + prod[524][5241] + prod[525][5251] + prod[526][5261] + prod[527][5271] + prod[528][5281] + prod[529][5291] + prod[530][5301] + prod[531][5311] + prod[532][5321] + prod[533][5331] + prod[534][5341] + prod[535][5351] + prod[536][5361] + prod[537][5371] + prod[538][5381] + prod[539][5391] + prod[540][5401] + prod[541][5411] + prod[542][5421] + prod[543][5431] + prod[544][5441] + prod[545][5451] + prod[546][5461] + prod[547][5471] + prod[548][5481] + prod[549][5491] + prod[550][5501] + prod[551][5511] + prod[552][5521] + prod[553][5531] + prod[554][5541] + prod[555][5551] + prod[556][5561] + prod[557][5571] + prod[558][5581] + prod[559][5591] + prod[560][5601] + prod[561][5611] + prod[562][5621] + prod[563][5631] + prod[564][5641] + prod[565][5651] + prod[566][5661] + prod[567][5671] + prod[568][5681] + prod[569][5691] + prod[570][5701] + prod[571][5711] + prod[572][5721] + prod[573][5731] + prod[574][5741] + prod[575][5751] + prod[576][5761] + prod[577][5771] + prod[578][5781] + prod[579][5791] + prod[580][5801] + prod[581][5811] + prod[582][5821] + prod[583][5831] + prod[584][5841] + prod[585][5851] + prod[586][5861] + prod[587][5871] + prod[588][5881] + prod[589][5891] + prod[590][5901] + prod[591][5911] + prod[592][5921] + prod[593][5931] + prod[594][5941] + prod[595][5951] + prod[596][5961] + prod[597][5971] + prod[598][5981] + prod[599][5991] + prod[600][6001] + prod[601][6011] + prod[602][6021] + prod[603][6031] + prod[604][6041] + prod[605][6051] + prod[606][6061] + prod[607][6071] + prod[608][6081] + prod[609][6091] + prod[610][6101] + prod[611][6111] + prod[612][6121] + prod[613][6131] + prod[614][6141] + prod[615][6151] + prod[616][6161] + prod[617][6171] + prod[618][6181] + prod[619][6191] + prod[620][6201] + prod[621][6211] + prod[622][6221] + prod[623][6231] + prod[624][6241] + prod[625][6251] + prod[626][6261] + prod[627][6271] + prod[628][6281] + prod[629][6291] + prod[630][6301] + prod[631][6311] + prod[632][6321] + prod[633][6331] + prod[634][6341] + prod[635][6351] + prod[636][6361] + prod[637][6371] + prod[638][6381] + prod[639][6391] + prod[640][6401] + prod[641][6411] + prod[642][6421] + prod[643][6431] + prod[644][6441] + prod[645][6451] + prod[646][6461] + prod[647][6471] + prod[648][6481] + prod[649][6491] + prod[650][6501] + prod[651][6511] + prod[652][6521] + prod[653][6531] + prod[654][6541] + prod[655][6551] + prod[656][6561] + prod[657][6571] + prod[658][6581] + prod[659][6591] + prod[660][6601] + prod[661][6611] + prod[662][6621] + prod[663][6631] + prod[664][6641] + prod[665][6651] + prod[666][6661] + prod[667][6671] + prod[668][6681] + prod[669][6691] + prod[670][6701] + prod[671][6711] + prod[672][6721] + prod[673][6731] + prod[674][6741] + prod[675][6751] + prod[676][6761] + prod[677][6771] + prod[678][6781] + prod[679][6791] + prod[680][6801] + prod[681][6811] + prod[682][6821] + prod[683][6831] + prod[684][6841] + prod[685][6851] + prod[686][6861] + prod[687][6871] + prod[688][6881] + prod[689][6891] + prod[690][6901] + prod[691][6911] + prod[692][6921] + prod[693][6931] + prod[694][6941] + prod[695][6951] + prod[696][6961] + prod[697][6971] + prod[698][6981] + prod[699][6991] + prod[700][7001] + prod[701][7011] + prod[702][7021] + prod[703][7031] + prod[704][7041] + prod[705][7051] + prod[706][7061] + prod[707][7071] + prod[708][7081] + prod[709][7091] + prod[710][7101] + prod[711][7111] + prod[712][7121] + prod[713][7131] + prod[714][7141] + prod[715][7151] + prod[716][7161] + prod[717][7171] + prod[718][7181] + prod[719][7191] + prod[720][7201] + prod[721][7211] + prod[722][7221] + prod[723][7231] + prod[724][7241] + prod[725][7251] + prod[726][7261] + prod[727][7271] + prod[728][7281] + prod[729][7291] + prod[730][7301] + prod[731][7311] + prod[732][7321] + prod[733][7331] + prod[734][7341] + prod[735][7351] + prod[736][7361] + prod[737][7371] + prod[738][7381] + prod[739][7391] + prod[740][7401] + prod[741][7411] + prod[742][7421] + prod[743][7431] + prod[744][7441] + prod[745][7451] + prod[746][7461] + prod[747][7471] + prod[748][7481] + prod[749][7491] + prod[750][7501] + prod[751][7511] + prod[752][7521] + prod[753][7531] + prod[754][7541] + prod[755][7551] + prod[756][7561] + prod[757][7571] + prod[758][7581] + prod[759][7591] + prod[760][7601] + prod[761][7611] + prod[762][7621] + prod[763][7631] + prod[764][7641] + prod[765][7651] + prod[766][7661] + prod[767][7671] + prod[768][7681] + prod[769][7691] + prod[770][7701] + prod[771][7711] + prod[772][7721] + prod[773][7731] + prod[774][7741] + prod[775][7751] + prod[776][7761] + prod[777][7771] + prod[778][7781] + prod[779][7791] + prod[780][7801] + prod[781][7811] + prod[782][7821] + prod[783][7831];
mul_temp[2] = prod[0][2] + prod[1][12] + prod[2][22] + prod[3][32] + prod[4][42] + prod[5][52] + prod[6][62] + prod[7][72] + prod[8][82] + prod[9][92] + prod[10][102] + prod[11][112] + prod[12][122] + prod[13][132] + prod[14][142] + prod[15][152] + prod[16][162] + prod[17][172] + prod[18][182] + prod[19][192] + prod[20][202] + prod[21][212] + prod[22][222] + prod[23][232] + prod[24][242] + prod[25][252] + prod[26][262] + prod[27][272] + prod[28][282] + prod[29][292] + prod[30][302] + prod[31][312] + prod[32][322] + prod[33][332] + prod[34][342] + prod[35][352] + prod[36][362] + prod[37][372] + prod[38][382] + prod[39][392] + prod[40][402] + prod[41][412] + prod[42][422] + prod[43][432] + prod[44][442] + prod[45][452] + prod[46][462] + prod[47][472] + prod[48][482] + prod[49][492] + prod[50][502] + prod[51][512] + prod[52][522] + prod[53][532] + prod[54][542] + prod[55][552] + prod[56][562] + prod[57][572] + prod[58][582] + prod[59][592] + prod[60][602] + prod[61][612] + prod[62][622] + prod[63][632] + prod[64][642] + prod[65][652] + prod[66][662] + prod[67][672] + prod[68][682] + prod[69][692] + prod[70][702] + prod[71][712] + prod[72][722] + prod[73][732] + prod[74][742] + prod[75][752] + prod[76][762] + prod[77][772] + prod[78][782] + prod[79][792] + prod[80][802] + prod[81][812] + prod[82][822] + prod[83][832] + prod[84][842] + prod[85][852] + prod[86][862] + prod[87][872] + prod[88][882] + prod[89][892] + prod[90][902] + prod[91][912] + prod[92][922] + prod[93][932] + prod[94][942] + prod[95][952] + prod[96][962] + prod[97][972] + prod[98][982] + prod[99][992] + prod[100][1002] + prod[101][1012] + prod[102][1022] + prod[103][1032] + prod[104][1042] + prod[105][1052] + prod[106][1062] + prod[107][1072] + prod[108][1082] + prod[109][1092] + prod[110][1102] + prod[111][1112] + prod[112][1122] + prod[113][1132] + prod[114][1142] + prod[115][1152] + prod[116][1162] + prod[117][1172] + prod[118][1182] + prod[119][1192] + prod[120][1202] + prod[121][1212] + prod[122][1222] + prod[123][1232] + prod[124][1242] + prod[125][1252] + prod[126][1262] + prod[127][1272] + prod[128][1282] + prod[129][1292] + prod[130][1302] + prod[131][1312] + prod[132][1322] + prod[133][1332] + prod[134][1342] + prod[135][1352] + prod[136][1362] + prod[137][1372] + prod[138][1382] + prod[139][1392] + prod[140][1402] + prod[141][1412] + prod[142][1422] + prod[143][1432] + prod[144][1442] + prod[145][1452] + prod[146][1462] + prod[147][1472] + prod[148][1482] + prod[149][1492] + prod[150][1502] + prod[151][1512] + prod[152][1522] + prod[153][1532] + prod[154][1542] + prod[155][1552] + prod[156][1562] + prod[157][1572] + prod[158][1582] + prod[159][1592] + prod[160][1602] + prod[161][1612] + prod[162][1622] + prod[163][1632] + prod[164][1642] + prod[165][1652] + prod[166][1662] + prod[167][1672] + prod[168][1682] + prod[169][1692] + prod[170][1702] + prod[171][1712] + prod[172][1722] + prod[173][1732] + prod[174][1742] + prod[175][1752] + prod[176][1762] + prod[177][1772] + prod[178][1782] + prod[179][1792] + prod[180][1802] + prod[181][1812] + prod[182][1822] + prod[183][1832] + prod[184][1842] + prod[185][1852] + prod[186][1862] + prod[187][1872] + prod[188][1882] + prod[189][1892] + prod[190][1902] + prod[191][1912] + prod[192][1922] + prod[193][1932] + prod[194][1942] + prod[195][1952] + prod[196][1962] + prod[197][1972] + prod[198][1982] + prod[199][1992] + prod[200][2002] + prod[201][2012] + prod[202][2022] + prod[203][2032] + prod[204][2042] + prod[205][2052] + prod[206][2062] + prod[207][2072] + prod[208][2082] + prod[209][2092] + prod[210][2102] + prod[211][2112] + prod[212][2122] + prod[213][2132] + prod[214][2142] + prod[215][2152] + prod[216][2162] + prod[217][2172] + prod[218][2182] + prod[219][2192] + prod[220][2202] + prod[221][2212] + prod[222][2222] + prod[223][2232] + prod[224][2242] + prod[225][2252] + prod[226][2262] + prod[227][2272] + prod[228][2282] + prod[229][2292] + prod[230][2302] + prod[231][2312] + prod[232][2322] + prod[233][2332] + prod[234][2342] + prod[235][2352] + prod[236][2362] + prod[237][2372] + prod[238][2382] + prod[239][2392] + prod[240][2402] + prod[241][2412] + prod[242][2422] + prod[243][2432] + prod[244][2442] + prod[245][2452] + prod[246][2462] + prod[247][2472] + prod[248][2482] + prod[249][2492] + prod[250][2502] + prod[251][2512] + prod[252][2522] + prod[253][2532] + prod[254][2542] + prod[255][2552] + prod[256][2562] + prod[257][2572] + prod[258][2582] + prod[259][2592] + prod[260][2602] + prod[261][2612] + prod[262][2622] + prod[263][2632] + prod[264][2642] + prod[265][2652] + prod[266][2662] + prod[267][2672] + prod[268][2682] + prod[269][2692] + prod[270][2702] + prod[271][2712] + prod[272][2722] + prod[273][2732] + prod[274][2742] + prod[275][2752] + prod[276][2762] + prod[277][2772] + prod[278][2782] + prod[279][2792] + prod[280][2802] + prod[281][2812] + prod[282][2822] + prod[283][2832] + prod[284][2842] + prod[285][2852] + prod[286][2862] + prod[287][2872] + prod[288][2882] + prod[289][2892] + prod[290][2902] + prod[291][2912] + prod[292][2922] + prod[293][2932] + prod[294][2942] + prod[295][2952] + prod[296][2962] + prod[297][2972] + prod[298][2982] + prod[299][2992] + prod[300][3002] + prod[301][3012] + prod[302][3022] + prod[303][3032] + prod[304][3042] + prod[305][3052] + prod[306][3062] + prod[307][3072] + prod[308][3082] + prod[309][3092] + prod[310][3102] + prod[311][3112] + prod[312][3122] + prod[313][3132] + prod[314][3142] + prod[315][3152] + prod[316][3162] + prod[317][3172] + prod[318][3182] + prod[319][3192] + prod[320][3202] + prod[321][3212] + prod[322][3222] + prod[323][3232] + prod[324][3242] + prod[325][3252] + prod[326][3262] + prod[327][3272] + prod[328][3282] + prod[329][3292] + prod[330][3302] + prod[331][3312] + prod[332][3322] + prod[333][3332] + prod[334][3342] + prod[335][3352] + prod[336][3362] + prod[337][3372] + prod[338][3382] + prod[339][3392] + prod[340][3402] + prod[341][3412] + prod[342][3422] + prod[343][3432] + prod[344][3442] + prod[345][3452] + prod[346][3462] + prod[347][3472] + prod[348][3482] + prod[349][3492] + prod[350][3502] + prod[351][3512] + prod[352][3522] + prod[353][3532] + prod[354][3542] + prod[355][3552] + prod[356][3562] + prod[357][3572] + prod[358][3582] + prod[359][3592] + prod[360][3602] + prod[361][3612] + prod[362][3622] + prod[363][3632] + prod[364][3642] + prod[365][3652] + prod[366][3662] + prod[367][3672] + prod[368][3682] + prod[369][3692] + prod[370][3702] + prod[371][3712] + prod[372][3722] + prod[373][3732] + prod[374][3742] + prod[375][3752] + prod[376][3762] + prod[377][3772] + prod[378][3782] + prod[379][3792] + prod[380][3802] + prod[381][3812] + prod[382][3822] + prod[383][3832] + prod[384][3842] + prod[385][3852] + prod[386][3862] + prod[387][3872] + prod[388][3882] + prod[389][3892] + prod[390][3902] + prod[391][3912] + prod[392][3922] + prod[393][3932] + prod[394][3942] + prod[395][3952] + prod[396][3962] + prod[397][3972] + prod[398][3982] + prod[399][3992] + prod[400][4002] + prod[401][4012] + prod[402][4022] + prod[403][4032] + prod[404][4042] + prod[405][4052] + prod[406][4062] + prod[407][4072] + prod[408][4082] + prod[409][4092] + prod[410][4102] + prod[411][4112] + prod[412][4122] + prod[413][4132] + prod[414][4142] + prod[415][4152] + prod[416][4162] + prod[417][4172] + prod[418][4182] + prod[419][4192] + prod[420][4202] + prod[421][4212] + prod[422][4222] + prod[423][4232] + prod[424][4242] + prod[425][4252] + prod[426][4262] + prod[427][4272] + prod[428][4282] + prod[429][4292] + prod[430][4302] + prod[431][4312] + prod[432][4322] + prod[433][4332] + prod[434][4342] + prod[435][4352] + prod[436][4362] + prod[437][4372] + prod[438][4382] + prod[439][4392] + prod[440][4402] + prod[441][4412] + prod[442][4422] + prod[443][4432] + prod[444][4442] + prod[445][4452] + prod[446][4462] + prod[447][4472] + prod[448][4482] + prod[449][4492] + prod[450][4502] + prod[451][4512] + prod[452][4522] + prod[453][4532] + prod[454][4542] + prod[455][4552] + prod[456][4562] + prod[457][4572] + prod[458][4582] + prod[459][4592] + prod[460][4602] + prod[461][4612] + prod[462][4622] + prod[463][4632] + prod[464][4642] + prod[465][4652] + prod[466][4662] + prod[467][4672] + prod[468][4682] + prod[469][4692] + prod[470][4702] + prod[471][4712] + prod[472][4722] + prod[473][4732] + prod[474][4742] + prod[475][4752] + prod[476][4762] + prod[477][4772] + prod[478][4782] + prod[479][4792] + prod[480][4802] + prod[481][4812] + prod[482][4822] + prod[483][4832] + prod[484][4842] + prod[485][4852] + prod[486][4862] + prod[487][4872] + prod[488][4882] + prod[489][4892] + prod[490][4902] + prod[491][4912] + prod[492][4922] + prod[493][4932] + prod[494][4942] + prod[495][4952] + prod[496][4962] + prod[497][4972] + prod[498][4982] + prod[499][4992] + prod[500][5002] + prod[501][5012] + prod[502][5022] + prod[503][5032] + prod[504][5042] + prod[505][5052] + prod[506][5062] + prod[507][5072] + prod[508][5082] + prod[509][5092] + prod[510][5102] + prod[511][5112] + prod[512][5122] + prod[513][5132] + prod[514][5142] + prod[515][5152] + prod[516][5162] + prod[517][5172] + prod[518][5182] + prod[519][5192] + prod[520][5202] + prod[521][5212] + prod[522][5222] + prod[523][5232] + prod[524][5242] + prod[525][5252] + prod[526][5262] + prod[527][5272] + prod[528][5282] + prod[529][5292] + prod[530][5302] + prod[531][5312] + prod[532][5322] + prod[533][5332] + prod[534][5342] + prod[535][5352] + prod[536][5362] + prod[537][5372] + prod[538][5382] + prod[539][5392] + prod[540][5402] + prod[541][5412] + prod[542][5422] + prod[543][5432] + prod[544][5442] + prod[545][5452] + prod[546][5462] + prod[547][5472] + prod[548][5482] + prod[549][5492] + prod[550][5502] + prod[551][5512] + prod[552][5522] + prod[553][5532] + prod[554][5542] + prod[555][5552] + prod[556][5562] + prod[557][5572] + prod[558][5582] + prod[559][5592] + prod[560][5602] + prod[561][5612] + prod[562][5622] + prod[563][5632] + prod[564][5642] + prod[565][5652] + prod[566][5662] + prod[567][5672] + prod[568][5682] + prod[569][5692] + prod[570][5702] + prod[571][5712] + prod[572][5722] + prod[573][5732] + prod[574][5742] + prod[575][5752] + prod[576][5762] + prod[577][5772] + prod[578][5782] + prod[579][5792] + prod[580][5802] + prod[581][5812] + prod[582][5822] + prod[583][5832] + prod[584][5842] + prod[585][5852] + prod[586][5862] + prod[587][5872] + prod[588][5882] + prod[589][5892] + prod[590][5902] + prod[591][5912] + prod[592][5922] + prod[593][5932] + prod[594][5942] + prod[595][5952] + prod[596][5962] + prod[597][5972] + prod[598][5982] + prod[599][5992] + prod[600][6002] + prod[601][6012] + prod[602][6022] + prod[603][6032] + prod[604][6042] + prod[605][6052] + prod[606][6062] + prod[607][6072] + prod[608][6082] + prod[609][6092] + prod[610][6102] + prod[611][6112] + prod[612][6122] + prod[613][6132] + prod[614][6142] + prod[615][6152] + prod[616][6162] + prod[617][6172] + prod[618][6182] + prod[619][6192] + prod[620][6202] + prod[621][6212] + prod[622][6222] + prod[623][6232] + prod[624][6242] + prod[625][6252] + prod[626][6262] + prod[627][6272] + prod[628][6282] + prod[629][6292] + prod[630][6302] + prod[631][6312] + prod[632][6322] + prod[633][6332] + prod[634][6342] + prod[635][6352] + prod[636][6362] + prod[637][6372] + prod[638][6382] + prod[639][6392] + prod[640][6402] + prod[641][6412] + prod[642][6422] + prod[643][6432] + prod[644][6442] + prod[645][6452] + prod[646][6462] + prod[647][6472] + prod[648][6482] + prod[649][6492] + prod[650][6502] + prod[651][6512] + prod[652][6522] + prod[653][6532] + prod[654][6542] + prod[655][6552] + prod[656][6562] + prod[657][6572] + prod[658][6582] + prod[659][6592] + prod[660][6602] + prod[661][6612] + prod[662][6622] + prod[663][6632] + prod[664][6642] + prod[665][6652] + prod[666][6662] + prod[667][6672] + prod[668][6682] + prod[669][6692] + prod[670][6702] + prod[671][6712] + prod[672][6722] + prod[673][6732] + prod[674][6742] + prod[675][6752] + prod[676][6762] + prod[677][6772] + prod[678][6782] + prod[679][6792] + prod[680][6802] + prod[681][6812] + prod[682][6822] + prod[683][6832] + prod[684][6842] + prod[685][6852] + prod[686][6862] + prod[687][6872] + prod[688][6882] + prod[689][6892] + prod[690][6902] + prod[691][6912] + prod[692][6922] + prod[693][6932] + prod[694][6942] + prod[695][6952] + prod[696][6962] + prod[697][6972] + prod[698][6982] + prod[699][6992] + prod[700][7002] + prod[701][7012] + prod[702][7022] + prod[703][7032] + prod[704][7042] + prod[705][7052] + prod[706][7062] + prod[707][7072] + prod[708][7082] + prod[709][7092] + prod[710][7102] + prod[711][7112] + prod[712][7122] + prod[713][7132] + prod[714][7142] + prod[715][7152] + prod[716][7162] + prod[717][7172] + prod[718][7182] + prod[719][7192] + prod[720][7202] + prod[721][7212] + prod[722][7222] + prod[723][7232] + prod[724][7242] + prod[725][7252] + prod[726][7262] + prod[727][7272] + prod[728][7282] + prod[729][7292] + prod[730][7302] + prod[731][7312] + prod[732][7322] + prod[733][7332] + prod[734][7342] + prod[735][7352] + prod[736][7362] + prod[737][7372] + prod[738][7382] + prod[739][7392] + prod[740][7402] + prod[741][7412] + prod[742][7422] + prod[743][7432] + prod[744][7442] + prod[745][7452] + prod[746][7462] + prod[747][7472] + prod[748][7482] + prod[749][7492] + prod[750][7502] + prod[751][7512] + prod[752][7522] + prod[753][7532] + prod[754][7542] + prod[755][7552] + prod[756][7562] + prod[757][7572] + prod[758][7582] + prod[759][7592] + prod[760][7602] + prod[761][7612] + prod[762][7622] + prod[763][7632] + prod[764][7642] + prod[765][7652] + prod[766][7662] + prod[767][7672] + prod[768][7682] + prod[769][7692] + prod[770][7702] + prod[771][7712] + prod[772][7722] + prod[773][7732] + prod[774][7742] + prod[775][7752] + prod[776][7762] + prod[777][7772] + prod[778][7782] + prod[779][7792] + prod[780][7802] + prod[781][7812] + prod[782][7822] + prod[783][7832];
mul_temp[3] = prod[0][3] + prod[1][13] + prod[2][23] + prod[3][33] + prod[4][43] + prod[5][53] + prod[6][63] + prod[7][73] + prod[8][83] + prod[9][93] + prod[10][103] + prod[11][113] + prod[12][123] + prod[13][133] + prod[14][143] + prod[15][153] + prod[16][163] + prod[17][173] + prod[18][183] + prod[19][193] + prod[20][203] + prod[21][213] + prod[22][223] + prod[23][233] + prod[24][243] + prod[25][253] + prod[26][263] + prod[27][273] + prod[28][283] + prod[29][293] + prod[30][303] + prod[31][313] + prod[32][323] + prod[33][333] + prod[34][343] + prod[35][353] + prod[36][363] + prod[37][373] + prod[38][383] + prod[39][393] + prod[40][403] + prod[41][413] + prod[42][423] + prod[43][433] + prod[44][443] + prod[45][453] + prod[46][463] + prod[47][473] + prod[48][483] + prod[49][493] + prod[50][503] + prod[51][513] + prod[52][523] + prod[53][533] + prod[54][543] + prod[55][553] + prod[56][563] + prod[57][573] + prod[58][583] + prod[59][593] + prod[60][603] + prod[61][613] + prod[62][623] + prod[63][633] + prod[64][643] + prod[65][653] + prod[66][663] + prod[67][673] + prod[68][683] + prod[69][693] + prod[70][703] + prod[71][713] + prod[72][723] + prod[73][733] + prod[74][743] + prod[75][753] + prod[76][763] + prod[77][773] + prod[78][783] + prod[79][793] + prod[80][803] + prod[81][813] + prod[82][823] + prod[83][833] + prod[84][843] + prod[85][853] + prod[86][863] + prod[87][873] + prod[88][883] + prod[89][893] + prod[90][903] + prod[91][913] + prod[92][923] + prod[93][933] + prod[94][943] + prod[95][953] + prod[96][963] + prod[97][973] + prod[98][983] + prod[99][993] + prod[100][1003] + prod[101][1013] + prod[102][1023] + prod[103][1033] + prod[104][1043] + prod[105][1053] + prod[106][1063] + prod[107][1073] + prod[108][1083] + prod[109][1093] + prod[110][1103] + prod[111][1113] + prod[112][1123] + prod[113][1133] + prod[114][1143] + prod[115][1153] + prod[116][1163] + prod[117][1173] + prod[118][1183] + prod[119][1193] + prod[120][1203] + prod[121][1213] + prod[122][1223] + prod[123][1233] + prod[124][1243] + prod[125][1253] + prod[126][1263] + prod[127][1273] + prod[128][1283] + prod[129][1293] + prod[130][1303] + prod[131][1313] + prod[132][1323] + prod[133][1333] + prod[134][1343] + prod[135][1353] + prod[136][1363] + prod[137][1373] + prod[138][1383] + prod[139][1393] + prod[140][1403] + prod[141][1413] + prod[142][1423] + prod[143][1433] + prod[144][1443] + prod[145][1453] + prod[146][1463] + prod[147][1473] + prod[148][1483] + prod[149][1493] + prod[150][1503] + prod[151][1513] + prod[152][1523] + prod[153][1533] + prod[154][1543] + prod[155][1553] + prod[156][1563] + prod[157][1573] + prod[158][1583] + prod[159][1593] + prod[160][1603] + prod[161][1613] + prod[162][1623] + prod[163][1633] + prod[164][1643] + prod[165][1653] + prod[166][1663] + prod[167][1673] + prod[168][1683] + prod[169][1693] + prod[170][1703] + prod[171][1713] + prod[172][1723] + prod[173][1733] + prod[174][1743] + prod[175][1753] + prod[176][1763] + prod[177][1773] + prod[178][1783] + prod[179][1793] + prod[180][1803] + prod[181][1813] + prod[182][1823] + prod[183][1833] + prod[184][1843] + prod[185][1853] + prod[186][1863] + prod[187][1873] + prod[188][1883] + prod[189][1893] + prod[190][1903] + prod[191][1913] + prod[192][1923] + prod[193][1933] + prod[194][1943] + prod[195][1953] + prod[196][1963] + prod[197][1973] + prod[198][1983] + prod[199][1993] + prod[200][2003] + prod[201][2013] + prod[202][2023] + prod[203][2033] + prod[204][2043] + prod[205][2053] + prod[206][2063] + prod[207][2073] + prod[208][2083] + prod[209][2093] + prod[210][2103] + prod[211][2113] + prod[212][2123] + prod[213][2133] + prod[214][2143] + prod[215][2153] + prod[216][2163] + prod[217][2173] + prod[218][2183] + prod[219][2193] + prod[220][2203] + prod[221][2213] + prod[222][2223] + prod[223][2233] + prod[224][2243] + prod[225][2253] + prod[226][2263] + prod[227][2273] + prod[228][2283] + prod[229][2293] + prod[230][2303] + prod[231][2313] + prod[232][2323] + prod[233][2333] + prod[234][2343] + prod[235][2353] + prod[236][2363] + prod[237][2373] + prod[238][2383] + prod[239][2393] + prod[240][2403] + prod[241][2413] + prod[242][2423] + prod[243][2433] + prod[244][2443] + prod[245][2453] + prod[246][2463] + prod[247][2473] + prod[248][2483] + prod[249][2493] + prod[250][2503] + prod[251][2513] + prod[252][2523] + prod[253][2533] + prod[254][2543] + prod[255][2553] + prod[256][2563] + prod[257][2573] + prod[258][2583] + prod[259][2593] + prod[260][2603] + prod[261][2613] + prod[262][2623] + prod[263][2633] + prod[264][2643] + prod[265][2653] + prod[266][2663] + prod[267][2673] + prod[268][2683] + prod[269][2693] + prod[270][2703] + prod[271][2713] + prod[272][2723] + prod[273][2733] + prod[274][2743] + prod[275][2753] + prod[276][2763] + prod[277][2773] + prod[278][2783] + prod[279][2793] + prod[280][2803] + prod[281][2813] + prod[282][2823] + prod[283][2833] + prod[284][2843] + prod[285][2853] + prod[286][2863] + prod[287][2873] + prod[288][2883] + prod[289][2893] + prod[290][2903] + prod[291][2913] + prod[292][2923] + prod[293][2933] + prod[294][2943] + prod[295][2953] + prod[296][2963] + prod[297][2973] + prod[298][2983] + prod[299][2993] + prod[300][3003] + prod[301][3013] + prod[302][3023] + prod[303][3033] + prod[304][3043] + prod[305][3053] + prod[306][3063] + prod[307][3073] + prod[308][3083] + prod[309][3093] + prod[310][3103] + prod[311][3113] + prod[312][3123] + prod[313][3133] + prod[314][3143] + prod[315][3153] + prod[316][3163] + prod[317][3173] + prod[318][3183] + prod[319][3193] + prod[320][3203] + prod[321][3213] + prod[322][3223] + prod[323][3233] + prod[324][3243] + prod[325][3253] + prod[326][3263] + prod[327][3273] + prod[328][3283] + prod[329][3293] + prod[330][3303] + prod[331][3313] + prod[332][3323] + prod[333][3333] + prod[334][3343] + prod[335][3353] + prod[336][3363] + prod[337][3373] + prod[338][3383] + prod[339][3393] + prod[340][3403] + prod[341][3413] + prod[342][3423] + prod[343][3433] + prod[344][3443] + prod[345][3453] + prod[346][3463] + prod[347][3473] + prod[348][3483] + prod[349][3493] + prod[350][3503] + prod[351][3513] + prod[352][3523] + prod[353][3533] + prod[354][3543] + prod[355][3553] + prod[356][3563] + prod[357][3573] + prod[358][3583] + prod[359][3593] + prod[360][3603] + prod[361][3613] + prod[362][3623] + prod[363][3633] + prod[364][3643] + prod[365][3653] + prod[366][3663] + prod[367][3673] + prod[368][3683] + prod[369][3693] + prod[370][3703] + prod[371][3713] + prod[372][3723] + prod[373][3733] + prod[374][3743] + prod[375][3753] + prod[376][3763] + prod[377][3773] + prod[378][3783] + prod[379][3793] + prod[380][3803] + prod[381][3813] + prod[382][3823] + prod[383][3833] + prod[384][3843] + prod[385][3853] + prod[386][3863] + prod[387][3873] + prod[388][3883] + prod[389][3893] + prod[390][3903] + prod[391][3913] + prod[392][3923] + prod[393][3933] + prod[394][3943] + prod[395][3953] + prod[396][3963] + prod[397][3973] + prod[398][3983] + prod[399][3993] + prod[400][4003] + prod[401][4013] + prod[402][4023] + prod[403][4033] + prod[404][4043] + prod[405][4053] + prod[406][4063] + prod[407][4073] + prod[408][4083] + prod[409][4093] + prod[410][4103] + prod[411][4113] + prod[412][4123] + prod[413][4133] + prod[414][4143] + prod[415][4153] + prod[416][4163] + prod[417][4173] + prod[418][4183] + prod[419][4193] + prod[420][4203] + prod[421][4213] + prod[422][4223] + prod[423][4233] + prod[424][4243] + prod[425][4253] + prod[426][4263] + prod[427][4273] + prod[428][4283] + prod[429][4293] + prod[430][4303] + prod[431][4313] + prod[432][4323] + prod[433][4333] + prod[434][4343] + prod[435][4353] + prod[436][4363] + prod[437][4373] + prod[438][4383] + prod[439][4393] + prod[440][4403] + prod[441][4413] + prod[442][4423] + prod[443][4433] + prod[444][4443] + prod[445][4453] + prod[446][4463] + prod[447][4473] + prod[448][4483] + prod[449][4493] + prod[450][4503] + prod[451][4513] + prod[452][4523] + prod[453][4533] + prod[454][4543] + prod[455][4553] + prod[456][4563] + prod[457][4573] + prod[458][4583] + prod[459][4593] + prod[460][4603] + prod[461][4613] + prod[462][4623] + prod[463][4633] + prod[464][4643] + prod[465][4653] + prod[466][4663] + prod[467][4673] + prod[468][4683] + prod[469][4693] + prod[470][4703] + prod[471][4713] + prod[472][4723] + prod[473][4733] + prod[474][4743] + prod[475][4753] + prod[476][4763] + prod[477][4773] + prod[478][4783] + prod[479][4793] + prod[480][4803] + prod[481][4813] + prod[482][4823] + prod[483][4833] + prod[484][4843] + prod[485][4853] + prod[486][4863] + prod[487][4873] + prod[488][4883] + prod[489][4893] + prod[490][4903] + prod[491][4913] + prod[492][4923] + prod[493][4933] + prod[494][4943] + prod[495][4953] + prod[496][4963] + prod[497][4973] + prod[498][4983] + prod[499][4993] + prod[500][5003] + prod[501][5013] + prod[502][5023] + prod[503][5033] + prod[504][5043] + prod[505][5053] + prod[506][5063] + prod[507][5073] + prod[508][5083] + prod[509][5093] + prod[510][5103] + prod[511][5113] + prod[512][5123] + prod[513][5133] + prod[514][5143] + prod[515][5153] + prod[516][5163] + prod[517][5173] + prod[518][5183] + prod[519][5193] + prod[520][5203] + prod[521][5213] + prod[522][5223] + prod[523][5233] + prod[524][5243] + prod[525][5253] + prod[526][5263] + prod[527][5273] + prod[528][5283] + prod[529][5293] + prod[530][5303] + prod[531][5313] + prod[532][5323] + prod[533][5333] + prod[534][5343] + prod[535][5353] + prod[536][5363] + prod[537][5373] + prod[538][5383] + prod[539][5393] + prod[540][5403] + prod[541][5413] + prod[542][5423] + prod[543][5433] + prod[544][5443] + prod[545][5453] + prod[546][5463] + prod[547][5473] + prod[548][5483] + prod[549][5493] + prod[550][5503] + prod[551][5513] + prod[552][5523] + prod[553][5533] + prod[554][5543] + prod[555][5553] + prod[556][5563] + prod[557][5573] + prod[558][5583] + prod[559][5593] + prod[560][5603] + prod[561][5613] + prod[562][5623] + prod[563][5633] + prod[564][5643] + prod[565][5653] + prod[566][5663] + prod[567][5673] + prod[568][5683] + prod[569][5693] + prod[570][5703] + prod[571][5713] + prod[572][5723] + prod[573][5733] + prod[574][5743] + prod[575][5753] + prod[576][5763] + prod[577][5773] + prod[578][5783] + prod[579][5793] + prod[580][5803] + prod[581][5813] + prod[582][5823] + prod[583][5833] + prod[584][5843] + prod[585][5853] + prod[586][5863] + prod[587][5873] + prod[588][5883] + prod[589][5893] + prod[590][5903] + prod[591][5913] + prod[592][5923] + prod[593][5933] + prod[594][5943] + prod[595][5953] + prod[596][5963] + prod[597][5973] + prod[598][5983] + prod[599][5993] + prod[600][6003] + prod[601][6013] + prod[602][6023] + prod[603][6033] + prod[604][6043] + prod[605][6053] + prod[606][6063] + prod[607][6073] + prod[608][6083] + prod[609][6093] + prod[610][6103] + prod[611][6113] + prod[612][6123] + prod[613][6133] + prod[614][6143] + prod[615][6153] + prod[616][6163] + prod[617][6173] + prod[618][6183] + prod[619][6193] + prod[620][6203] + prod[621][6213] + prod[622][6223] + prod[623][6233] + prod[624][6243] + prod[625][6253] + prod[626][6263] + prod[627][6273] + prod[628][6283] + prod[629][6293] + prod[630][6303] + prod[631][6313] + prod[632][6323] + prod[633][6333] + prod[634][6343] + prod[635][6353] + prod[636][6363] + prod[637][6373] + prod[638][6383] + prod[639][6393] + prod[640][6403] + prod[641][6413] + prod[642][6423] + prod[643][6433] + prod[644][6443] + prod[645][6453] + prod[646][6463] + prod[647][6473] + prod[648][6483] + prod[649][6493] + prod[650][6503] + prod[651][6513] + prod[652][6523] + prod[653][6533] + prod[654][6543] + prod[655][6553] + prod[656][6563] + prod[657][6573] + prod[658][6583] + prod[659][6593] + prod[660][6603] + prod[661][6613] + prod[662][6623] + prod[663][6633] + prod[664][6643] + prod[665][6653] + prod[666][6663] + prod[667][6673] + prod[668][6683] + prod[669][6693] + prod[670][6703] + prod[671][6713] + prod[672][6723] + prod[673][6733] + prod[674][6743] + prod[675][6753] + prod[676][6763] + prod[677][6773] + prod[678][6783] + prod[679][6793] + prod[680][6803] + prod[681][6813] + prod[682][6823] + prod[683][6833] + prod[684][6843] + prod[685][6853] + prod[686][6863] + prod[687][6873] + prod[688][6883] + prod[689][6893] + prod[690][6903] + prod[691][6913] + prod[692][6923] + prod[693][6933] + prod[694][6943] + prod[695][6953] + prod[696][6963] + prod[697][6973] + prod[698][6983] + prod[699][6993] + prod[700][7003] + prod[701][7013] + prod[702][7023] + prod[703][7033] + prod[704][7043] + prod[705][7053] + prod[706][7063] + prod[707][7073] + prod[708][7083] + prod[709][7093] + prod[710][7103] + prod[711][7113] + prod[712][7123] + prod[713][7133] + prod[714][7143] + prod[715][7153] + prod[716][7163] + prod[717][7173] + prod[718][7183] + prod[719][7193] + prod[720][7203] + prod[721][7213] + prod[722][7223] + prod[723][7233] + prod[724][7243] + prod[725][7253] + prod[726][7263] + prod[727][7273] + prod[728][7283] + prod[729][7293] + prod[730][7303] + prod[731][7313] + prod[732][7323] + prod[733][7333] + prod[734][7343] + prod[735][7353] + prod[736][7363] + prod[737][7373] + prod[738][7383] + prod[739][7393] + prod[740][7403] + prod[741][7413] + prod[742][7423] + prod[743][7433] + prod[744][7443] + prod[745][7453] + prod[746][7463] + prod[747][7473] + prod[748][7483] + prod[749][7493] + prod[750][7503] + prod[751][7513] + prod[752][7523] + prod[753][7533] + prod[754][7543] + prod[755][7553] + prod[756][7563] + prod[757][7573] + prod[758][7583] + prod[759][7593] + prod[760][7603] + prod[761][7613] + prod[762][7623] + prod[763][7633] + prod[764][7643] + prod[765][7653] + prod[766][7663] + prod[767][7673] + prod[768][7683] + prod[769][7693] + prod[770][7703] + prod[771][7713] + prod[772][7723] + prod[773][7733] + prod[774][7743] + prod[775][7753] + prod[776][7763] + prod[777][7773] + prod[778][7783] + prod[779][7793] + prod[780][7803] + prod[781][7813] + prod[782][7823] + prod[783][7833];
mul_temp[4] = prod[0][4] + prod[1][14] + prod[2][24] + prod[3][34] + prod[4][44] + prod[5][54] + prod[6][64] + prod[7][74] + prod[8][84] + prod[9][94] + prod[10][104] + prod[11][114] + prod[12][124] + prod[13][134] + prod[14][144] + prod[15][154] + prod[16][164] + prod[17][174] + prod[18][184] + prod[19][194] + prod[20][204] + prod[21][214] + prod[22][224] + prod[23][234] + prod[24][244] + prod[25][254] + prod[26][264] + prod[27][274] + prod[28][284] + prod[29][294] + prod[30][304] + prod[31][314] + prod[32][324] + prod[33][334] + prod[34][344] + prod[35][354] + prod[36][364] + prod[37][374] + prod[38][384] + prod[39][394] + prod[40][404] + prod[41][414] + prod[42][424] + prod[43][434] + prod[44][444] + prod[45][454] + prod[46][464] + prod[47][474] + prod[48][484] + prod[49][494] + prod[50][504] + prod[51][514] + prod[52][524] + prod[53][534] + prod[54][544] + prod[55][554] + prod[56][564] + prod[57][574] + prod[58][584] + prod[59][594] + prod[60][604] + prod[61][614] + prod[62][624] + prod[63][634] + prod[64][644] + prod[65][654] + prod[66][664] + prod[67][674] + prod[68][684] + prod[69][694] + prod[70][704] + prod[71][714] + prod[72][724] + prod[73][734] + prod[74][744] + prod[75][754] + prod[76][764] + prod[77][774] + prod[78][784] + prod[79][794] + prod[80][804] + prod[81][814] + prod[82][824] + prod[83][834] + prod[84][844] + prod[85][854] + prod[86][864] + prod[87][874] + prod[88][884] + prod[89][894] + prod[90][904] + prod[91][914] + prod[92][924] + prod[93][934] + prod[94][944] + prod[95][954] + prod[96][964] + prod[97][974] + prod[98][984] + prod[99][994] + prod[100][1004] + prod[101][1014] + prod[102][1024] + prod[103][1034] + prod[104][1044] + prod[105][1054] + prod[106][1064] + prod[107][1074] + prod[108][1084] + prod[109][1094] + prod[110][1104] + prod[111][1114] + prod[112][1124] + prod[113][1134] + prod[114][1144] + prod[115][1154] + prod[116][1164] + prod[117][1174] + prod[118][1184] + prod[119][1194] + prod[120][1204] + prod[121][1214] + prod[122][1224] + prod[123][1234] + prod[124][1244] + prod[125][1254] + prod[126][1264] + prod[127][1274] + prod[128][1284] + prod[129][1294] + prod[130][1304] + prod[131][1314] + prod[132][1324] + prod[133][1334] + prod[134][1344] + prod[135][1354] + prod[136][1364] + prod[137][1374] + prod[138][1384] + prod[139][1394] + prod[140][1404] + prod[141][1414] + prod[142][1424] + prod[143][1434] + prod[144][1444] + prod[145][1454] + prod[146][1464] + prod[147][1474] + prod[148][1484] + prod[149][1494] + prod[150][1504] + prod[151][1514] + prod[152][1524] + prod[153][1534] + prod[154][1544] + prod[155][1554] + prod[156][1564] + prod[157][1574] + prod[158][1584] + prod[159][1594] + prod[160][1604] + prod[161][1614] + prod[162][1624] + prod[163][1634] + prod[164][1644] + prod[165][1654] + prod[166][1664] + prod[167][1674] + prod[168][1684] + prod[169][1694] + prod[170][1704] + prod[171][1714] + prod[172][1724] + prod[173][1734] + prod[174][1744] + prod[175][1754] + prod[176][1764] + prod[177][1774] + prod[178][1784] + prod[179][1794] + prod[180][1804] + prod[181][1814] + prod[182][1824] + prod[183][1834] + prod[184][1844] + prod[185][1854] + prod[186][1864] + prod[187][1874] + prod[188][1884] + prod[189][1894] + prod[190][1904] + prod[191][1914] + prod[192][1924] + prod[193][1934] + prod[194][1944] + prod[195][1954] + prod[196][1964] + prod[197][1974] + prod[198][1984] + prod[199][1994] + prod[200][2004] + prod[201][2014] + prod[202][2024] + prod[203][2034] + prod[204][2044] + prod[205][2054] + prod[206][2064] + prod[207][2074] + prod[208][2084] + prod[209][2094] + prod[210][2104] + prod[211][2114] + prod[212][2124] + prod[213][2134] + prod[214][2144] + prod[215][2154] + prod[216][2164] + prod[217][2174] + prod[218][2184] + prod[219][2194] + prod[220][2204] + prod[221][2214] + prod[222][2224] + prod[223][2234] + prod[224][2244] + prod[225][2254] + prod[226][2264] + prod[227][2274] + prod[228][2284] + prod[229][2294] + prod[230][2304] + prod[231][2314] + prod[232][2324] + prod[233][2334] + prod[234][2344] + prod[235][2354] + prod[236][2364] + prod[237][2374] + prod[238][2384] + prod[239][2394] + prod[240][2404] + prod[241][2414] + prod[242][2424] + prod[243][2434] + prod[244][2444] + prod[245][2454] + prod[246][2464] + prod[247][2474] + prod[248][2484] + prod[249][2494] + prod[250][2504] + prod[251][2514] + prod[252][2524] + prod[253][2534] + prod[254][2544] + prod[255][2554] + prod[256][2564] + prod[257][2574] + prod[258][2584] + prod[259][2594] + prod[260][2604] + prod[261][2614] + prod[262][2624] + prod[263][2634] + prod[264][2644] + prod[265][2654] + prod[266][2664] + prod[267][2674] + prod[268][2684] + prod[269][2694] + prod[270][2704] + prod[271][2714] + prod[272][2724] + prod[273][2734] + prod[274][2744] + prod[275][2754] + prod[276][2764] + prod[277][2774] + prod[278][2784] + prod[279][2794] + prod[280][2804] + prod[281][2814] + prod[282][2824] + prod[283][2834] + prod[284][2844] + prod[285][2854] + prod[286][2864] + prod[287][2874] + prod[288][2884] + prod[289][2894] + prod[290][2904] + prod[291][2914] + prod[292][2924] + prod[293][2934] + prod[294][2944] + prod[295][2954] + prod[296][2964] + prod[297][2974] + prod[298][2984] + prod[299][2994] + prod[300][3004] + prod[301][3014] + prod[302][3024] + prod[303][3034] + prod[304][3044] + prod[305][3054] + prod[306][3064] + prod[307][3074] + prod[308][3084] + prod[309][3094] + prod[310][3104] + prod[311][3114] + prod[312][3124] + prod[313][3134] + prod[314][3144] + prod[315][3154] + prod[316][3164] + prod[317][3174] + prod[318][3184] + prod[319][3194] + prod[320][3204] + prod[321][3214] + prod[322][3224] + prod[323][3234] + prod[324][3244] + prod[325][3254] + prod[326][3264] + prod[327][3274] + prod[328][3284] + prod[329][3294] + prod[330][3304] + prod[331][3314] + prod[332][3324] + prod[333][3334] + prod[334][3344] + prod[335][3354] + prod[336][3364] + prod[337][3374] + prod[338][3384] + prod[339][3394] + prod[340][3404] + prod[341][3414] + prod[342][3424] + prod[343][3434] + prod[344][3444] + prod[345][3454] + prod[346][3464] + prod[347][3474] + prod[348][3484] + prod[349][3494] + prod[350][3504] + prod[351][3514] + prod[352][3524] + prod[353][3534] + prod[354][3544] + prod[355][3554] + prod[356][3564] + prod[357][3574] + prod[358][3584] + prod[359][3594] + prod[360][3604] + prod[361][3614] + prod[362][3624] + prod[363][3634] + prod[364][3644] + prod[365][3654] + prod[366][3664] + prod[367][3674] + prod[368][3684] + prod[369][3694] + prod[370][3704] + prod[371][3714] + prod[372][3724] + prod[373][3734] + prod[374][3744] + prod[375][3754] + prod[376][3764] + prod[377][3774] + prod[378][3784] + prod[379][3794] + prod[380][3804] + prod[381][3814] + prod[382][3824] + prod[383][3834] + prod[384][3844] + prod[385][3854] + prod[386][3864] + prod[387][3874] + prod[388][3884] + prod[389][3894] + prod[390][3904] + prod[391][3914] + prod[392][3924] + prod[393][3934] + prod[394][3944] + prod[395][3954] + prod[396][3964] + prod[397][3974] + prod[398][3984] + prod[399][3994] + prod[400][4004] + prod[401][4014] + prod[402][4024] + prod[403][4034] + prod[404][4044] + prod[405][4054] + prod[406][4064] + prod[407][4074] + prod[408][4084] + prod[409][4094] + prod[410][4104] + prod[411][4114] + prod[412][4124] + prod[413][4134] + prod[414][4144] + prod[415][4154] + prod[416][4164] + prod[417][4174] + prod[418][4184] + prod[419][4194] + prod[420][4204] + prod[421][4214] + prod[422][4224] + prod[423][4234] + prod[424][4244] + prod[425][4254] + prod[426][4264] + prod[427][4274] + prod[428][4284] + prod[429][4294] + prod[430][4304] + prod[431][4314] + prod[432][4324] + prod[433][4334] + prod[434][4344] + prod[435][4354] + prod[436][4364] + prod[437][4374] + prod[438][4384] + prod[439][4394] + prod[440][4404] + prod[441][4414] + prod[442][4424] + prod[443][4434] + prod[444][4444] + prod[445][4454] + prod[446][4464] + prod[447][4474] + prod[448][4484] + prod[449][4494] + prod[450][4504] + prod[451][4514] + prod[452][4524] + prod[453][4534] + prod[454][4544] + prod[455][4554] + prod[456][4564] + prod[457][4574] + prod[458][4584] + prod[459][4594] + prod[460][4604] + prod[461][4614] + prod[462][4624] + prod[463][4634] + prod[464][4644] + prod[465][4654] + prod[466][4664] + prod[467][4674] + prod[468][4684] + prod[469][4694] + prod[470][4704] + prod[471][4714] + prod[472][4724] + prod[473][4734] + prod[474][4744] + prod[475][4754] + prod[476][4764] + prod[477][4774] + prod[478][4784] + prod[479][4794] + prod[480][4804] + prod[481][4814] + prod[482][4824] + prod[483][4834] + prod[484][4844] + prod[485][4854] + prod[486][4864] + prod[487][4874] + prod[488][4884] + prod[489][4894] + prod[490][4904] + prod[491][4914] + prod[492][4924] + prod[493][4934] + prod[494][4944] + prod[495][4954] + prod[496][4964] + prod[497][4974] + prod[498][4984] + prod[499][4994] + prod[500][5004] + prod[501][5014] + prod[502][5024] + prod[503][5034] + prod[504][5044] + prod[505][5054] + prod[506][5064] + prod[507][5074] + prod[508][5084] + prod[509][5094] + prod[510][5104] + prod[511][5114] + prod[512][5124] + prod[513][5134] + prod[514][5144] + prod[515][5154] + prod[516][5164] + prod[517][5174] + prod[518][5184] + prod[519][5194] + prod[520][5204] + prod[521][5214] + prod[522][5224] + prod[523][5234] + prod[524][5244] + prod[525][5254] + prod[526][5264] + prod[527][5274] + prod[528][5284] + prod[529][5294] + prod[530][5304] + prod[531][5314] + prod[532][5324] + prod[533][5334] + prod[534][5344] + prod[535][5354] + prod[536][5364] + prod[537][5374] + prod[538][5384] + prod[539][5394] + prod[540][5404] + prod[541][5414] + prod[542][5424] + prod[543][5434] + prod[544][5444] + prod[545][5454] + prod[546][5464] + prod[547][5474] + prod[548][5484] + prod[549][5494] + prod[550][5504] + prod[551][5514] + prod[552][5524] + prod[553][5534] + prod[554][5544] + prod[555][5554] + prod[556][5564] + prod[557][5574] + prod[558][5584] + prod[559][5594] + prod[560][5604] + prod[561][5614] + prod[562][5624] + prod[563][5634] + prod[564][5644] + prod[565][5654] + prod[566][5664] + prod[567][5674] + prod[568][5684] + prod[569][5694] + prod[570][5704] + prod[571][5714] + prod[572][5724] + prod[573][5734] + prod[574][5744] + prod[575][5754] + prod[576][5764] + prod[577][5774] + prod[578][5784] + prod[579][5794] + prod[580][5804] + prod[581][5814] + prod[582][5824] + prod[583][5834] + prod[584][5844] + prod[585][5854] + prod[586][5864] + prod[587][5874] + prod[588][5884] + prod[589][5894] + prod[590][5904] + prod[591][5914] + prod[592][5924] + prod[593][5934] + prod[594][5944] + prod[595][5954] + prod[596][5964] + prod[597][5974] + prod[598][5984] + prod[599][5994] + prod[600][6004] + prod[601][6014] + prod[602][6024] + prod[603][6034] + prod[604][6044] + prod[605][6054] + prod[606][6064] + prod[607][6074] + prod[608][6084] + prod[609][6094] + prod[610][6104] + prod[611][6114] + prod[612][6124] + prod[613][6134] + prod[614][6144] + prod[615][6154] + prod[616][6164] + prod[617][6174] + prod[618][6184] + prod[619][6194] + prod[620][6204] + prod[621][6214] + prod[622][6224] + prod[623][6234] + prod[624][6244] + prod[625][6254] + prod[626][6264] + prod[627][6274] + prod[628][6284] + prod[629][6294] + prod[630][6304] + prod[631][6314] + prod[632][6324] + prod[633][6334] + prod[634][6344] + prod[635][6354] + prod[636][6364] + prod[637][6374] + prod[638][6384] + prod[639][6394] + prod[640][6404] + prod[641][6414] + prod[642][6424] + prod[643][6434] + prod[644][6444] + prod[645][6454] + prod[646][6464] + prod[647][6474] + prod[648][6484] + prod[649][6494] + prod[650][6504] + prod[651][6514] + prod[652][6524] + prod[653][6534] + prod[654][6544] + prod[655][6554] + prod[656][6564] + prod[657][6574] + prod[658][6584] + prod[659][6594] + prod[660][6604] + prod[661][6614] + prod[662][6624] + prod[663][6634] + prod[664][6644] + prod[665][6654] + prod[666][6664] + prod[667][6674] + prod[668][6684] + prod[669][6694] + prod[670][6704] + prod[671][6714] + prod[672][6724] + prod[673][6734] + prod[674][6744] + prod[675][6754] + prod[676][6764] + prod[677][6774] + prod[678][6784] + prod[679][6794] + prod[680][6804] + prod[681][6814] + prod[682][6824] + prod[683][6834] + prod[684][6844] + prod[685][6854] + prod[686][6864] + prod[687][6874] + prod[688][6884] + prod[689][6894] + prod[690][6904] + prod[691][6914] + prod[692][6924] + prod[693][6934] + prod[694][6944] + prod[695][6954] + prod[696][6964] + prod[697][6974] + prod[698][6984] + prod[699][6994] + prod[700][7004] + prod[701][7014] + prod[702][7024] + prod[703][7034] + prod[704][7044] + prod[705][7054] + prod[706][7064] + prod[707][7074] + prod[708][7084] + prod[709][7094] + prod[710][7104] + prod[711][7114] + prod[712][7124] + prod[713][7134] + prod[714][7144] + prod[715][7154] + prod[716][7164] + prod[717][7174] + prod[718][7184] + prod[719][7194] + prod[720][7204] + prod[721][7214] + prod[722][7224] + prod[723][7234] + prod[724][7244] + prod[725][7254] + prod[726][7264] + prod[727][7274] + prod[728][7284] + prod[729][7294] + prod[730][7304] + prod[731][7314] + prod[732][7324] + prod[733][7334] + prod[734][7344] + prod[735][7354] + prod[736][7364] + prod[737][7374] + prod[738][7384] + prod[739][7394] + prod[740][7404] + prod[741][7414] + prod[742][7424] + prod[743][7434] + prod[744][7444] + prod[745][7454] + prod[746][7464] + prod[747][7474] + prod[748][7484] + prod[749][7494] + prod[750][7504] + prod[751][7514] + prod[752][7524] + prod[753][7534] + prod[754][7544] + prod[755][7554] + prod[756][7564] + prod[757][7574] + prod[758][7584] + prod[759][7594] + prod[760][7604] + prod[761][7614] + prod[762][7624] + prod[763][7634] + prod[764][7644] + prod[765][7654] + prod[766][7664] + prod[767][7674] + prod[768][7684] + prod[769][7694] + prod[770][7704] + prod[771][7714] + prod[772][7724] + prod[773][7734] + prod[774][7744] + prod[775][7754] + prod[776][7764] + prod[777][7774] + prod[778][7784] + prod[779][7794] + prod[780][7804] + prod[781][7814] + prod[782][7824] + prod[783][7834];
mul_temp[5] = prod[0][5] + prod[1][15] + prod[2][25] + prod[3][35] + prod[4][45] + prod[5][55] + prod[6][65] + prod[7][75] + prod[8][85] + prod[9][95] + prod[10][105] + prod[11][115] + prod[12][125] + prod[13][135] + prod[14][145] + prod[15][155] + prod[16][165] + prod[17][175] + prod[18][185] + prod[19][195] + prod[20][205] + prod[21][215] + prod[22][225] + prod[23][235] + prod[24][245] + prod[25][255] + prod[26][265] + prod[27][275] + prod[28][285] + prod[29][295] + prod[30][305] + prod[31][315] + prod[32][325] + prod[33][335] + prod[34][345] + prod[35][355] + prod[36][365] + prod[37][375] + prod[38][385] + prod[39][395] + prod[40][405] + prod[41][415] + prod[42][425] + prod[43][435] + prod[44][445] + prod[45][455] + prod[46][465] + prod[47][475] + prod[48][485] + prod[49][495] + prod[50][505] + prod[51][515] + prod[52][525] + prod[53][535] + prod[54][545] + prod[55][555] + prod[56][565] + prod[57][575] + prod[58][585] + prod[59][595] + prod[60][605] + prod[61][615] + prod[62][625] + prod[63][635] + prod[64][645] + prod[65][655] + prod[66][665] + prod[67][675] + prod[68][685] + prod[69][695] + prod[70][705] + prod[71][715] + prod[72][725] + prod[73][735] + prod[74][745] + prod[75][755] + prod[76][765] + prod[77][775] + prod[78][785] + prod[79][795] + prod[80][805] + prod[81][815] + prod[82][825] + prod[83][835] + prod[84][845] + prod[85][855] + prod[86][865] + prod[87][875] + prod[88][885] + prod[89][895] + prod[90][905] + prod[91][915] + prod[92][925] + prod[93][935] + prod[94][945] + prod[95][955] + prod[96][965] + prod[97][975] + prod[98][985] + prod[99][995] + prod[100][1005] + prod[101][1015] + prod[102][1025] + prod[103][1035] + prod[104][1045] + prod[105][1055] + prod[106][1065] + prod[107][1075] + prod[108][1085] + prod[109][1095] + prod[110][1105] + prod[111][1115] + prod[112][1125] + prod[113][1135] + prod[114][1145] + prod[115][1155] + prod[116][1165] + prod[117][1175] + prod[118][1185] + prod[119][1195] + prod[120][1205] + prod[121][1215] + prod[122][1225] + prod[123][1235] + prod[124][1245] + prod[125][1255] + prod[126][1265] + prod[127][1275] + prod[128][1285] + prod[129][1295] + prod[130][1305] + prod[131][1315] + prod[132][1325] + prod[133][1335] + prod[134][1345] + prod[135][1355] + prod[136][1365] + prod[137][1375] + prod[138][1385] + prod[139][1395] + prod[140][1405] + prod[141][1415] + prod[142][1425] + prod[143][1435] + prod[144][1445] + prod[145][1455] + prod[146][1465] + prod[147][1475] + prod[148][1485] + prod[149][1495] + prod[150][1505] + prod[151][1515] + prod[152][1525] + prod[153][1535] + prod[154][1545] + prod[155][1555] + prod[156][1565] + prod[157][1575] + prod[158][1585] + prod[159][1595] + prod[160][1605] + prod[161][1615] + prod[162][1625] + prod[163][1635] + prod[164][1645] + prod[165][1655] + prod[166][1665] + prod[167][1675] + prod[168][1685] + prod[169][1695] + prod[170][1705] + prod[171][1715] + prod[172][1725] + prod[173][1735] + prod[174][1745] + prod[175][1755] + prod[176][1765] + prod[177][1775] + prod[178][1785] + prod[179][1795] + prod[180][1805] + prod[181][1815] + prod[182][1825] + prod[183][1835] + prod[184][1845] + prod[185][1855] + prod[186][1865] + prod[187][1875] + prod[188][1885] + prod[189][1895] + prod[190][1905] + prod[191][1915] + prod[192][1925] + prod[193][1935] + prod[194][1945] + prod[195][1955] + prod[196][1965] + prod[197][1975] + prod[198][1985] + prod[199][1995] + prod[200][2005] + prod[201][2015] + prod[202][2025] + prod[203][2035] + prod[204][2045] + prod[205][2055] + prod[206][2065] + prod[207][2075] + prod[208][2085] + prod[209][2095] + prod[210][2105] + prod[211][2115] + prod[212][2125] + prod[213][2135] + prod[214][2145] + prod[215][2155] + prod[216][2165] + prod[217][2175] + prod[218][2185] + prod[219][2195] + prod[220][2205] + prod[221][2215] + prod[222][2225] + prod[223][2235] + prod[224][2245] + prod[225][2255] + prod[226][2265] + prod[227][2275] + prod[228][2285] + prod[229][2295] + prod[230][2305] + prod[231][2315] + prod[232][2325] + prod[233][2335] + prod[234][2345] + prod[235][2355] + prod[236][2365] + prod[237][2375] + prod[238][2385] + prod[239][2395] + prod[240][2405] + prod[241][2415] + prod[242][2425] + prod[243][2435] + prod[244][2445] + prod[245][2455] + prod[246][2465] + prod[247][2475] + prod[248][2485] + prod[249][2495] + prod[250][2505] + prod[251][2515] + prod[252][2525] + prod[253][2535] + prod[254][2545] + prod[255][2555] + prod[256][2565] + prod[257][2575] + prod[258][2585] + prod[259][2595] + prod[260][2605] + prod[261][2615] + prod[262][2625] + prod[263][2635] + prod[264][2645] + prod[265][2655] + prod[266][2665] + prod[267][2675] + prod[268][2685] + prod[269][2695] + prod[270][2705] + prod[271][2715] + prod[272][2725] + prod[273][2735] + prod[274][2745] + prod[275][2755] + prod[276][2765] + prod[277][2775] + prod[278][2785] + prod[279][2795] + prod[280][2805] + prod[281][2815] + prod[282][2825] + prod[283][2835] + prod[284][2845] + prod[285][2855] + prod[286][2865] + prod[287][2875] + prod[288][2885] + prod[289][2895] + prod[290][2905] + prod[291][2915] + prod[292][2925] + prod[293][2935] + prod[294][2945] + prod[295][2955] + prod[296][2965] + prod[297][2975] + prod[298][2985] + prod[299][2995] + prod[300][3005] + prod[301][3015] + prod[302][3025] + prod[303][3035] + prod[304][3045] + prod[305][3055] + prod[306][3065] + prod[307][3075] + prod[308][3085] + prod[309][3095] + prod[310][3105] + prod[311][3115] + prod[312][3125] + prod[313][3135] + prod[314][3145] + prod[315][3155] + prod[316][3165] + prod[317][3175] + prod[318][3185] + prod[319][3195] + prod[320][3205] + prod[321][3215] + prod[322][3225] + prod[323][3235] + prod[324][3245] + prod[325][3255] + prod[326][3265] + prod[327][3275] + prod[328][3285] + prod[329][3295] + prod[330][3305] + prod[331][3315] + prod[332][3325] + prod[333][3335] + prod[334][3345] + prod[335][3355] + prod[336][3365] + prod[337][3375] + prod[338][3385] + prod[339][3395] + prod[340][3405] + prod[341][3415] + prod[342][3425] + prod[343][3435] + prod[344][3445] + prod[345][3455] + prod[346][3465] + prod[347][3475] + prod[348][3485] + prod[349][3495] + prod[350][3505] + prod[351][3515] + prod[352][3525] + prod[353][3535] + prod[354][3545] + prod[355][3555] + prod[356][3565] + prod[357][3575] + prod[358][3585] + prod[359][3595] + prod[360][3605] + prod[361][3615] + prod[362][3625] + prod[363][3635] + prod[364][3645] + prod[365][3655] + prod[366][3665] + prod[367][3675] + prod[368][3685] + prod[369][3695] + prod[370][3705] + prod[371][3715] + prod[372][3725] + prod[373][3735] + prod[374][3745] + prod[375][3755] + prod[376][3765] + prod[377][3775] + prod[378][3785] + prod[379][3795] + prod[380][3805] + prod[381][3815] + prod[382][3825] + prod[383][3835] + prod[384][3845] + prod[385][3855] + prod[386][3865] + prod[387][3875] + prod[388][3885] + prod[389][3895] + prod[390][3905] + prod[391][3915] + prod[392][3925] + prod[393][3935] + prod[394][3945] + prod[395][3955] + prod[396][3965] + prod[397][3975] + prod[398][3985] + prod[399][3995] + prod[400][4005] + prod[401][4015] + prod[402][4025] + prod[403][4035] + prod[404][4045] + prod[405][4055] + prod[406][4065] + prod[407][4075] + prod[408][4085] + prod[409][4095] + prod[410][4105] + prod[411][4115] + prod[412][4125] + prod[413][4135] + prod[414][4145] + prod[415][4155] + prod[416][4165] + prod[417][4175] + prod[418][4185] + prod[419][4195] + prod[420][4205] + prod[421][4215] + prod[422][4225] + prod[423][4235] + prod[424][4245] + prod[425][4255] + prod[426][4265] + prod[427][4275] + prod[428][4285] + prod[429][4295] + prod[430][4305] + prod[431][4315] + prod[432][4325] + prod[433][4335] + prod[434][4345] + prod[435][4355] + prod[436][4365] + prod[437][4375] + prod[438][4385] + prod[439][4395] + prod[440][4405] + prod[441][4415] + prod[442][4425] + prod[443][4435] + prod[444][4445] + prod[445][4455] + prod[446][4465] + prod[447][4475] + prod[448][4485] + prod[449][4495] + prod[450][4505] + prod[451][4515] + prod[452][4525] + prod[453][4535] + prod[454][4545] + prod[455][4555] + prod[456][4565] + prod[457][4575] + prod[458][4585] + prod[459][4595] + prod[460][4605] + prod[461][4615] + prod[462][4625] + prod[463][4635] + prod[464][4645] + prod[465][4655] + prod[466][4665] + prod[467][4675] + prod[468][4685] + prod[469][4695] + prod[470][4705] + prod[471][4715] + prod[472][4725] + prod[473][4735] + prod[474][4745] + prod[475][4755] + prod[476][4765] + prod[477][4775] + prod[478][4785] + prod[479][4795] + prod[480][4805] + prod[481][4815] + prod[482][4825] + prod[483][4835] + prod[484][4845] + prod[485][4855] + prod[486][4865] + prod[487][4875] + prod[488][4885] + prod[489][4895] + prod[490][4905] + prod[491][4915] + prod[492][4925] + prod[493][4935] + prod[494][4945] + prod[495][4955] + prod[496][4965] + prod[497][4975] + prod[498][4985] + prod[499][4995] + prod[500][5005] + prod[501][5015] + prod[502][5025] + prod[503][5035] + prod[504][5045] + prod[505][5055] + prod[506][5065] + prod[507][5075] + prod[508][5085] + prod[509][5095] + prod[510][5105] + prod[511][5115] + prod[512][5125] + prod[513][5135] + prod[514][5145] + prod[515][5155] + prod[516][5165] + prod[517][5175] + prod[518][5185] + prod[519][5195] + prod[520][5205] + prod[521][5215] + prod[522][5225] + prod[523][5235] + prod[524][5245] + prod[525][5255] + prod[526][5265] + prod[527][5275] + prod[528][5285] + prod[529][5295] + prod[530][5305] + prod[531][5315] + prod[532][5325] + prod[533][5335] + prod[534][5345] + prod[535][5355] + prod[536][5365] + prod[537][5375] + prod[538][5385] + prod[539][5395] + prod[540][5405] + prod[541][5415] + prod[542][5425] + prod[543][5435] + prod[544][5445] + prod[545][5455] + prod[546][5465] + prod[547][5475] + prod[548][5485] + prod[549][5495] + prod[550][5505] + prod[551][5515] + prod[552][5525] + prod[553][5535] + prod[554][5545] + prod[555][5555] + prod[556][5565] + prod[557][5575] + prod[558][5585] + prod[559][5595] + prod[560][5605] + prod[561][5615] + prod[562][5625] + prod[563][5635] + prod[564][5645] + prod[565][5655] + prod[566][5665] + prod[567][5675] + prod[568][5685] + prod[569][5695] + prod[570][5705] + prod[571][5715] + prod[572][5725] + prod[573][5735] + prod[574][5745] + prod[575][5755] + prod[576][5765] + prod[577][5775] + prod[578][5785] + prod[579][5795] + prod[580][5805] + prod[581][5815] + prod[582][5825] + prod[583][5835] + prod[584][5845] + prod[585][5855] + prod[586][5865] + prod[587][5875] + prod[588][5885] + prod[589][5895] + prod[590][5905] + prod[591][5915] + prod[592][5925] + prod[593][5935] + prod[594][5945] + prod[595][5955] + prod[596][5965] + prod[597][5975] + prod[598][5985] + prod[599][5995] + prod[600][6005] + prod[601][6015] + prod[602][6025] + prod[603][6035] + prod[604][6045] + prod[605][6055] + prod[606][6065] + prod[607][6075] + prod[608][6085] + prod[609][6095] + prod[610][6105] + prod[611][6115] + prod[612][6125] + prod[613][6135] + prod[614][6145] + prod[615][6155] + prod[616][6165] + prod[617][6175] + prod[618][6185] + prod[619][6195] + prod[620][6205] + prod[621][6215] + prod[622][6225] + prod[623][6235] + prod[624][6245] + prod[625][6255] + prod[626][6265] + prod[627][6275] + prod[628][6285] + prod[629][6295] + prod[630][6305] + prod[631][6315] + prod[632][6325] + prod[633][6335] + prod[634][6345] + prod[635][6355] + prod[636][6365] + prod[637][6375] + prod[638][6385] + prod[639][6395] + prod[640][6405] + prod[641][6415] + prod[642][6425] + prod[643][6435] + prod[644][6445] + prod[645][6455] + prod[646][6465] + prod[647][6475] + prod[648][6485] + prod[649][6495] + prod[650][6505] + prod[651][6515] + prod[652][6525] + prod[653][6535] + prod[654][6545] + prod[655][6555] + prod[656][6565] + prod[657][6575] + prod[658][6585] + prod[659][6595] + prod[660][6605] + prod[661][6615] + prod[662][6625] + prod[663][6635] + prod[664][6645] + prod[665][6655] + prod[666][6665] + prod[667][6675] + prod[668][6685] + prod[669][6695] + prod[670][6705] + prod[671][6715] + prod[672][6725] + prod[673][6735] + prod[674][6745] + prod[675][6755] + prod[676][6765] + prod[677][6775] + prod[678][6785] + prod[679][6795] + prod[680][6805] + prod[681][6815] + prod[682][6825] + prod[683][6835] + prod[684][6845] + prod[685][6855] + prod[686][6865] + prod[687][6875] + prod[688][6885] + prod[689][6895] + prod[690][6905] + prod[691][6915] + prod[692][6925] + prod[693][6935] + prod[694][6945] + prod[695][6955] + prod[696][6965] + prod[697][6975] + prod[698][6985] + prod[699][6995] + prod[700][7005] + prod[701][7015] + prod[702][7025] + prod[703][7035] + prod[704][7045] + prod[705][7055] + prod[706][7065] + prod[707][7075] + prod[708][7085] + prod[709][7095] + prod[710][7105] + prod[711][7115] + prod[712][7125] + prod[713][7135] + prod[714][7145] + prod[715][7155] + prod[716][7165] + prod[717][7175] + prod[718][7185] + prod[719][7195] + prod[720][7205] + prod[721][7215] + prod[722][7225] + prod[723][7235] + prod[724][7245] + prod[725][7255] + prod[726][7265] + prod[727][7275] + prod[728][7285] + prod[729][7295] + prod[730][7305] + prod[731][7315] + prod[732][7325] + prod[733][7335] + prod[734][7345] + prod[735][7355] + prod[736][7365] + prod[737][7375] + prod[738][7385] + prod[739][7395] + prod[740][7405] + prod[741][7415] + prod[742][7425] + prod[743][7435] + prod[744][7445] + prod[745][7455] + prod[746][7465] + prod[747][7475] + prod[748][7485] + prod[749][7495] + prod[750][7505] + prod[751][7515] + prod[752][7525] + prod[753][7535] + prod[754][7545] + prod[755][7555] + prod[756][7565] + prod[757][7575] + prod[758][7585] + prod[759][7595] + prod[760][7605] + prod[761][7615] + prod[762][7625] + prod[763][7635] + prod[764][7645] + prod[765][7655] + prod[766][7665] + prod[767][7675] + prod[768][7685] + prod[769][7695] + prod[770][7705] + prod[771][7715] + prod[772][7725] + prod[773][7735] + prod[774][7745] + prod[775][7755] + prod[776][7765] + prod[777][7775] + prod[778][7785] + prod[779][7795] + prod[780][7805] + prod[781][7815] + prod[782][7825] + prod[783][7835];
mul_temp[6] = prod[0][6] + prod[1][16] + prod[2][26] + prod[3][36] + prod[4][46] + prod[5][56] + prod[6][66] + prod[7][76] + prod[8][86] + prod[9][96] + prod[10][106] + prod[11][116] + prod[12][126] + prod[13][136] + prod[14][146] + prod[15][156] + prod[16][166] + prod[17][176] + prod[18][186] + prod[19][196] + prod[20][206] + prod[21][216] + prod[22][226] + prod[23][236] + prod[24][246] + prod[25][256] + prod[26][266] + prod[27][276] + prod[28][286] + prod[29][296] + prod[30][306] + prod[31][316] + prod[32][326] + prod[33][336] + prod[34][346] + prod[35][356] + prod[36][366] + prod[37][376] + prod[38][386] + prod[39][396] + prod[40][406] + prod[41][416] + prod[42][426] + prod[43][436] + prod[44][446] + prod[45][456] + prod[46][466] + prod[47][476] + prod[48][486] + prod[49][496] + prod[50][506] + prod[51][516] + prod[52][526] + prod[53][536] + prod[54][546] + prod[55][556] + prod[56][566] + prod[57][576] + prod[58][586] + prod[59][596] + prod[60][606] + prod[61][616] + prod[62][626] + prod[63][636] + prod[64][646] + prod[65][656] + prod[66][666] + prod[67][676] + prod[68][686] + prod[69][696] + prod[70][706] + prod[71][716] + prod[72][726] + prod[73][736] + prod[74][746] + prod[75][756] + prod[76][766] + prod[77][776] + prod[78][786] + prod[79][796] + prod[80][806] + prod[81][816] + prod[82][826] + prod[83][836] + prod[84][846] + prod[85][856] + prod[86][866] + prod[87][876] + prod[88][886] + prod[89][896] + prod[90][906] + prod[91][916] + prod[92][926] + prod[93][936] + prod[94][946] + prod[95][956] + prod[96][966] + prod[97][976] + prod[98][986] + prod[99][996] + prod[100][1006] + prod[101][1016] + prod[102][1026] + prod[103][1036] + prod[104][1046] + prod[105][1056] + prod[106][1066] + prod[107][1076] + prod[108][1086] + prod[109][1096] + prod[110][1106] + prod[111][1116] + prod[112][1126] + prod[113][1136] + prod[114][1146] + prod[115][1156] + prod[116][1166] + prod[117][1176] + prod[118][1186] + prod[119][1196] + prod[120][1206] + prod[121][1216] + prod[122][1226] + prod[123][1236] + prod[124][1246] + prod[125][1256] + prod[126][1266] + prod[127][1276] + prod[128][1286] + prod[129][1296] + prod[130][1306] + prod[131][1316] + prod[132][1326] + prod[133][1336] + prod[134][1346] + prod[135][1356] + prod[136][1366] + prod[137][1376] + prod[138][1386] + prod[139][1396] + prod[140][1406] + prod[141][1416] + prod[142][1426] + prod[143][1436] + prod[144][1446] + prod[145][1456] + prod[146][1466] + prod[147][1476] + prod[148][1486] + prod[149][1496] + prod[150][1506] + prod[151][1516] + prod[152][1526] + prod[153][1536] + prod[154][1546] + prod[155][1556] + prod[156][1566] + prod[157][1576] + prod[158][1586] + prod[159][1596] + prod[160][1606] + prod[161][1616] + prod[162][1626] + prod[163][1636] + prod[164][1646] + prod[165][1656] + prod[166][1666] + prod[167][1676] + prod[168][1686] + prod[169][1696] + prod[170][1706] + prod[171][1716] + prod[172][1726] + prod[173][1736] + prod[174][1746] + prod[175][1756] + prod[176][1766] + prod[177][1776] + prod[178][1786] + prod[179][1796] + prod[180][1806] + prod[181][1816] + prod[182][1826] + prod[183][1836] + prod[184][1846] + prod[185][1856] + prod[186][1866] + prod[187][1876] + prod[188][1886] + prod[189][1896] + prod[190][1906] + prod[191][1916] + prod[192][1926] + prod[193][1936] + prod[194][1946] + prod[195][1956] + prod[196][1966] + prod[197][1976] + prod[198][1986] + prod[199][1996] + prod[200][2006] + prod[201][2016] + prod[202][2026] + prod[203][2036] + prod[204][2046] + prod[205][2056] + prod[206][2066] + prod[207][2076] + prod[208][2086] + prod[209][2096] + prod[210][2106] + prod[211][2116] + prod[212][2126] + prod[213][2136] + prod[214][2146] + prod[215][2156] + prod[216][2166] + prod[217][2176] + prod[218][2186] + prod[219][2196] + prod[220][2206] + prod[221][2216] + prod[222][2226] + prod[223][2236] + prod[224][2246] + prod[225][2256] + prod[226][2266] + prod[227][2276] + prod[228][2286] + prod[229][2296] + prod[230][2306] + prod[231][2316] + prod[232][2326] + prod[233][2336] + prod[234][2346] + prod[235][2356] + prod[236][2366] + prod[237][2376] + prod[238][2386] + prod[239][2396] + prod[240][2406] + prod[241][2416] + prod[242][2426] + prod[243][2436] + prod[244][2446] + prod[245][2456] + prod[246][2466] + prod[247][2476] + prod[248][2486] + prod[249][2496] + prod[250][2506] + prod[251][2516] + prod[252][2526] + prod[253][2536] + prod[254][2546] + prod[255][2556] + prod[256][2566] + prod[257][2576] + prod[258][2586] + prod[259][2596] + prod[260][2606] + prod[261][2616] + prod[262][2626] + prod[263][2636] + prod[264][2646] + prod[265][2656] + prod[266][2666] + prod[267][2676] + prod[268][2686] + prod[269][2696] + prod[270][2706] + prod[271][2716] + prod[272][2726] + prod[273][2736] + prod[274][2746] + prod[275][2756] + prod[276][2766] + prod[277][2776] + prod[278][2786] + prod[279][2796] + prod[280][2806] + prod[281][2816] + prod[282][2826] + prod[283][2836] + prod[284][2846] + prod[285][2856] + prod[286][2866] + prod[287][2876] + prod[288][2886] + prod[289][2896] + prod[290][2906] + prod[291][2916] + prod[292][2926] + prod[293][2936] + prod[294][2946] + prod[295][2956] + prod[296][2966] + prod[297][2976] + prod[298][2986] + prod[299][2996] + prod[300][3006] + prod[301][3016] + prod[302][3026] + prod[303][3036] + prod[304][3046] + prod[305][3056] + prod[306][3066] + prod[307][3076] + prod[308][3086] + prod[309][3096] + prod[310][3106] + prod[311][3116] + prod[312][3126] + prod[313][3136] + prod[314][3146] + prod[315][3156] + prod[316][3166] + prod[317][3176] + prod[318][3186] + prod[319][3196] + prod[320][3206] + prod[321][3216] + prod[322][3226] + prod[323][3236] + prod[324][3246] + prod[325][3256] + prod[326][3266] + prod[327][3276] + prod[328][3286] + prod[329][3296] + prod[330][3306] + prod[331][3316] + prod[332][3326] + prod[333][3336] + prod[334][3346] + prod[335][3356] + prod[336][3366] + prod[337][3376] + prod[338][3386] + prod[339][3396] + prod[340][3406] + prod[341][3416] + prod[342][3426] + prod[343][3436] + prod[344][3446] + prod[345][3456] + prod[346][3466] + prod[347][3476] + prod[348][3486] + prod[349][3496] + prod[350][3506] + prod[351][3516] + prod[352][3526] + prod[353][3536] + prod[354][3546] + prod[355][3556] + prod[356][3566] + prod[357][3576] + prod[358][3586] + prod[359][3596] + prod[360][3606] + prod[361][3616] + prod[362][3626] + prod[363][3636] + prod[364][3646] + prod[365][3656] + prod[366][3666] + prod[367][3676] + prod[368][3686] + prod[369][3696] + prod[370][3706] + prod[371][3716] + prod[372][3726] + prod[373][3736] + prod[374][3746] + prod[375][3756] + prod[376][3766] + prod[377][3776] + prod[378][3786] + prod[379][3796] + prod[380][3806] + prod[381][3816] + prod[382][3826] + prod[383][3836] + prod[384][3846] + prod[385][3856] + prod[386][3866] + prod[387][3876] + prod[388][3886] + prod[389][3896] + prod[390][3906] + prod[391][3916] + prod[392][3926] + prod[393][3936] + prod[394][3946] + prod[395][3956] + prod[396][3966] + prod[397][3976] + prod[398][3986] + prod[399][3996] + prod[400][4006] + prod[401][4016] + prod[402][4026] + prod[403][4036] + prod[404][4046] + prod[405][4056] + prod[406][4066] + prod[407][4076] + prod[408][4086] + prod[409][4096] + prod[410][4106] + prod[411][4116] + prod[412][4126] + prod[413][4136] + prod[414][4146] + prod[415][4156] + prod[416][4166] + prod[417][4176] + prod[418][4186] + prod[419][4196] + prod[420][4206] + prod[421][4216] + prod[422][4226] + prod[423][4236] + prod[424][4246] + prod[425][4256] + prod[426][4266] + prod[427][4276] + prod[428][4286] + prod[429][4296] + prod[430][4306] + prod[431][4316] + prod[432][4326] + prod[433][4336] + prod[434][4346] + prod[435][4356] + prod[436][4366] + prod[437][4376] + prod[438][4386] + prod[439][4396] + prod[440][4406] + prod[441][4416] + prod[442][4426] + prod[443][4436] + prod[444][4446] + prod[445][4456] + prod[446][4466] + prod[447][4476] + prod[448][4486] + prod[449][4496] + prod[450][4506] + prod[451][4516] + prod[452][4526] + prod[453][4536] + prod[454][4546] + prod[455][4556] + prod[456][4566] + prod[457][4576] + prod[458][4586] + prod[459][4596] + prod[460][4606] + prod[461][4616] + prod[462][4626] + prod[463][4636] + prod[464][4646] + prod[465][4656] + prod[466][4666] + prod[467][4676] + prod[468][4686] + prod[469][4696] + prod[470][4706] + prod[471][4716] + prod[472][4726] + prod[473][4736] + prod[474][4746] + prod[475][4756] + prod[476][4766] + prod[477][4776] + prod[478][4786] + prod[479][4796] + prod[480][4806] + prod[481][4816] + prod[482][4826] + prod[483][4836] + prod[484][4846] + prod[485][4856] + prod[486][4866] + prod[487][4876] + prod[488][4886] + prod[489][4896] + prod[490][4906] + prod[491][4916] + prod[492][4926] + prod[493][4936] + prod[494][4946] + prod[495][4956] + prod[496][4966] + prod[497][4976] + prod[498][4986] + prod[499][4996] + prod[500][5006] + prod[501][5016] + prod[502][5026] + prod[503][5036] + prod[504][5046] + prod[505][5056] + prod[506][5066] + prod[507][5076] + prod[508][5086] + prod[509][5096] + prod[510][5106] + prod[511][5116] + prod[512][5126] + prod[513][5136] + prod[514][5146] + prod[515][5156] + prod[516][5166] + prod[517][5176] + prod[518][5186] + prod[519][5196] + prod[520][5206] + prod[521][5216] + prod[522][5226] + prod[523][5236] + prod[524][5246] + prod[525][5256] + prod[526][5266] + prod[527][5276] + prod[528][5286] + prod[529][5296] + prod[530][5306] + prod[531][5316] + prod[532][5326] + prod[533][5336] + prod[534][5346] + prod[535][5356] + prod[536][5366] + prod[537][5376] + prod[538][5386] + prod[539][5396] + prod[540][5406] + prod[541][5416] + prod[542][5426] + prod[543][5436] + prod[544][5446] + prod[545][5456] + prod[546][5466] + prod[547][5476] + prod[548][5486] + prod[549][5496] + prod[550][5506] + prod[551][5516] + prod[552][5526] + prod[553][5536] + prod[554][5546] + prod[555][5556] + prod[556][5566] + prod[557][5576] + prod[558][5586] + prod[559][5596] + prod[560][5606] + prod[561][5616] + prod[562][5626] + prod[563][5636] + prod[564][5646] + prod[565][5656] + prod[566][5666] + prod[567][5676] + prod[568][5686] + prod[569][5696] + prod[570][5706] + prod[571][5716] + prod[572][5726] + prod[573][5736] + prod[574][5746] + prod[575][5756] + prod[576][5766] + prod[577][5776] + prod[578][5786] + prod[579][5796] + prod[580][5806] + prod[581][5816] + prod[582][5826] + prod[583][5836] + prod[584][5846] + prod[585][5856] + prod[586][5866] + prod[587][5876] + prod[588][5886] + prod[589][5896] + prod[590][5906] + prod[591][5916] + prod[592][5926] + prod[593][5936] + prod[594][5946] + prod[595][5956] + prod[596][5966] + prod[597][5976] + prod[598][5986] + prod[599][5996] + prod[600][6006] + prod[601][6016] + prod[602][6026] + prod[603][6036] + prod[604][6046] + prod[605][6056] + prod[606][6066] + prod[607][6076] + prod[608][6086] + prod[609][6096] + prod[610][6106] + prod[611][6116] + prod[612][6126] + prod[613][6136] + prod[614][6146] + prod[615][6156] + prod[616][6166] + prod[617][6176] + prod[618][6186] + prod[619][6196] + prod[620][6206] + prod[621][6216] + prod[622][6226] + prod[623][6236] + prod[624][6246] + prod[625][6256] + prod[626][6266] + prod[627][6276] + prod[628][6286] + prod[629][6296] + prod[630][6306] + prod[631][6316] + prod[632][6326] + prod[633][6336] + prod[634][6346] + prod[635][6356] + prod[636][6366] + prod[637][6376] + prod[638][6386] + prod[639][6396] + prod[640][6406] + prod[641][6416] + prod[642][6426] + prod[643][6436] + prod[644][6446] + prod[645][6456] + prod[646][6466] + prod[647][6476] + prod[648][6486] + prod[649][6496] + prod[650][6506] + prod[651][6516] + prod[652][6526] + prod[653][6536] + prod[654][6546] + prod[655][6556] + prod[656][6566] + prod[657][6576] + prod[658][6586] + prod[659][6596] + prod[660][6606] + prod[661][6616] + prod[662][6626] + prod[663][6636] + prod[664][6646] + prod[665][6656] + prod[666][6666] + prod[667][6676] + prod[668][6686] + prod[669][6696] + prod[670][6706] + prod[671][6716] + prod[672][6726] + prod[673][6736] + prod[674][6746] + prod[675][6756] + prod[676][6766] + prod[677][6776] + prod[678][6786] + prod[679][6796] + prod[680][6806] + prod[681][6816] + prod[682][6826] + prod[683][6836] + prod[684][6846] + prod[685][6856] + prod[686][6866] + prod[687][6876] + prod[688][6886] + prod[689][6896] + prod[690][6906] + prod[691][6916] + prod[692][6926] + prod[693][6936] + prod[694][6946] + prod[695][6956] + prod[696][6966] + prod[697][6976] + prod[698][6986] + prod[699][6996] + prod[700][7006] + prod[701][7016] + prod[702][7026] + prod[703][7036] + prod[704][7046] + prod[705][7056] + prod[706][7066] + prod[707][7076] + prod[708][7086] + prod[709][7096] + prod[710][7106] + prod[711][7116] + prod[712][7126] + prod[713][7136] + prod[714][7146] + prod[715][7156] + prod[716][7166] + prod[717][7176] + prod[718][7186] + prod[719][7196] + prod[720][7206] + prod[721][7216] + prod[722][7226] + prod[723][7236] + prod[724][7246] + prod[725][7256] + prod[726][7266] + prod[727][7276] + prod[728][7286] + prod[729][7296] + prod[730][7306] + prod[731][7316] + prod[732][7326] + prod[733][7336] + prod[734][7346] + prod[735][7356] + prod[736][7366] + prod[737][7376] + prod[738][7386] + prod[739][7396] + prod[740][7406] + prod[741][7416] + prod[742][7426] + prod[743][7436] + prod[744][7446] + prod[745][7456] + prod[746][7466] + prod[747][7476] + prod[748][7486] + prod[749][7496] + prod[750][7506] + prod[751][7516] + prod[752][7526] + prod[753][7536] + prod[754][7546] + prod[755][7556] + prod[756][7566] + prod[757][7576] + prod[758][7586] + prod[759][7596] + prod[760][7606] + prod[761][7616] + prod[762][7626] + prod[763][7636] + prod[764][7646] + prod[765][7656] + prod[766][7666] + prod[767][7676] + prod[768][7686] + prod[769][7696] + prod[770][7706] + prod[771][7716] + prod[772][7726] + prod[773][7736] + prod[774][7746] + prod[775][7756] + prod[776][7766] + prod[777][7776] + prod[778][7786] + prod[779][7796] + prod[780][7806] + prod[781][7816] + prod[782][7826] + prod[783][7836];
mul_temp[7] = prod[0][7] + prod[1][17] + prod[2][27] + prod[3][37] + prod[4][47] + prod[5][57] + prod[6][67] + prod[7][77] + prod[8][87] + prod[9][97] + prod[10][107] + prod[11][117] + prod[12][127] + prod[13][137] + prod[14][147] + prod[15][157] + prod[16][167] + prod[17][177] + prod[18][187] + prod[19][197] + prod[20][207] + prod[21][217] + prod[22][227] + prod[23][237] + prod[24][247] + prod[25][257] + prod[26][267] + prod[27][277] + prod[28][287] + prod[29][297] + prod[30][307] + prod[31][317] + prod[32][327] + prod[33][337] + prod[34][347] + prod[35][357] + prod[36][367] + prod[37][377] + prod[38][387] + prod[39][397] + prod[40][407] + prod[41][417] + prod[42][427] + prod[43][437] + prod[44][447] + prod[45][457] + prod[46][467] + prod[47][477] + prod[48][487] + prod[49][497] + prod[50][507] + prod[51][517] + prod[52][527] + prod[53][537] + prod[54][547] + prod[55][557] + prod[56][567] + prod[57][577] + prod[58][587] + prod[59][597] + prod[60][607] + prod[61][617] + prod[62][627] + prod[63][637] + prod[64][647] + prod[65][657] + prod[66][667] + prod[67][677] + prod[68][687] + prod[69][697] + prod[70][707] + prod[71][717] + prod[72][727] + prod[73][737] + prod[74][747] + prod[75][757] + prod[76][767] + prod[77][777] + prod[78][787] + prod[79][797] + prod[80][807] + prod[81][817] + prod[82][827] + prod[83][837] + prod[84][847] + prod[85][857] + prod[86][867] + prod[87][877] + prod[88][887] + prod[89][897] + prod[90][907] + prod[91][917] + prod[92][927] + prod[93][937] + prod[94][947] + prod[95][957] + prod[96][967] + prod[97][977] + prod[98][987] + prod[99][997] + prod[100][1007] + prod[101][1017] + prod[102][1027] + prod[103][1037] + prod[104][1047] + prod[105][1057] + prod[106][1067] + prod[107][1077] + prod[108][1087] + prod[109][1097] + prod[110][1107] + prod[111][1117] + prod[112][1127] + prod[113][1137] + prod[114][1147] + prod[115][1157] + prod[116][1167] + prod[117][1177] + prod[118][1187] + prod[119][1197] + prod[120][1207] + prod[121][1217] + prod[122][1227] + prod[123][1237] + prod[124][1247] + prod[125][1257] + prod[126][1267] + prod[127][1277] + prod[128][1287] + prod[129][1297] + prod[130][1307] + prod[131][1317] + prod[132][1327] + prod[133][1337] + prod[134][1347] + prod[135][1357] + prod[136][1367] + prod[137][1377] + prod[138][1387] + prod[139][1397] + prod[140][1407] + prod[141][1417] + prod[142][1427] + prod[143][1437] + prod[144][1447] + prod[145][1457] + prod[146][1467] + prod[147][1477] + prod[148][1487] + prod[149][1497] + prod[150][1507] + prod[151][1517] + prod[152][1527] + prod[153][1537] + prod[154][1547] + prod[155][1557] + prod[156][1567] + prod[157][1577] + prod[158][1587] + prod[159][1597] + prod[160][1607] + prod[161][1617] + prod[162][1627] + prod[163][1637] + prod[164][1647] + prod[165][1657] + prod[166][1667] + prod[167][1677] + prod[168][1687] + prod[169][1697] + prod[170][1707] + prod[171][1717] + prod[172][1727] + prod[173][1737] + prod[174][1747] + prod[175][1757] + prod[176][1767] + prod[177][1777] + prod[178][1787] + prod[179][1797] + prod[180][1807] + prod[181][1817] + prod[182][1827] + prod[183][1837] + prod[184][1847] + prod[185][1857] + prod[186][1867] + prod[187][1877] + prod[188][1887] + prod[189][1897] + prod[190][1907] + prod[191][1917] + prod[192][1927] + prod[193][1937] + prod[194][1947] + prod[195][1957] + prod[196][1967] + prod[197][1977] + prod[198][1987] + prod[199][1997] + prod[200][2007] + prod[201][2017] + prod[202][2027] + prod[203][2037] + prod[204][2047] + prod[205][2057] + prod[206][2067] + prod[207][2077] + prod[208][2087] + prod[209][2097] + prod[210][2107] + prod[211][2117] + prod[212][2127] + prod[213][2137] + prod[214][2147] + prod[215][2157] + prod[216][2167] + prod[217][2177] + prod[218][2187] + prod[219][2197] + prod[220][2207] + prod[221][2217] + prod[222][2227] + prod[223][2237] + prod[224][2247] + prod[225][2257] + prod[226][2267] + prod[227][2277] + prod[228][2287] + prod[229][2297] + prod[230][2307] + prod[231][2317] + prod[232][2327] + prod[233][2337] + prod[234][2347] + prod[235][2357] + prod[236][2367] + prod[237][2377] + prod[238][2387] + prod[239][2397] + prod[240][2407] + prod[241][2417] + prod[242][2427] + prod[243][2437] + prod[244][2447] + prod[245][2457] + prod[246][2467] + prod[247][2477] + prod[248][2487] + prod[249][2497] + prod[250][2507] + prod[251][2517] + prod[252][2527] + prod[253][2537] + prod[254][2547] + prod[255][2557] + prod[256][2567] + prod[257][2577] + prod[258][2587] + prod[259][2597] + prod[260][2607] + prod[261][2617] + prod[262][2627] + prod[263][2637] + prod[264][2647] + prod[265][2657] + prod[266][2667] + prod[267][2677] + prod[268][2687] + prod[269][2697] + prod[270][2707] + prod[271][2717] + prod[272][2727] + prod[273][2737] + prod[274][2747] + prod[275][2757] + prod[276][2767] + prod[277][2777] + prod[278][2787] + prod[279][2797] + prod[280][2807] + prod[281][2817] + prod[282][2827] + prod[283][2837] + prod[284][2847] + prod[285][2857] + prod[286][2867] + prod[287][2877] + prod[288][2887] + prod[289][2897] + prod[290][2907] + prod[291][2917] + prod[292][2927] + prod[293][2937] + prod[294][2947] + prod[295][2957] + prod[296][2967] + prod[297][2977] + prod[298][2987] + prod[299][2997] + prod[300][3007] + prod[301][3017] + prod[302][3027] + prod[303][3037] + prod[304][3047] + prod[305][3057] + prod[306][3067] + prod[307][3077] + prod[308][3087] + prod[309][3097] + prod[310][3107] + prod[311][3117] + prod[312][3127] + prod[313][3137] + prod[314][3147] + prod[315][3157] + prod[316][3167] + prod[317][3177] + prod[318][3187] + prod[319][3197] + prod[320][3207] + prod[321][3217] + prod[322][3227] + prod[323][3237] + prod[324][3247] + prod[325][3257] + prod[326][3267] + prod[327][3277] + prod[328][3287] + prod[329][3297] + prod[330][3307] + prod[331][3317] + prod[332][3327] + prod[333][3337] + prod[334][3347] + prod[335][3357] + prod[336][3367] + prod[337][3377] + prod[338][3387] + prod[339][3397] + prod[340][3407] + prod[341][3417] + prod[342][3427] + prod[343][3437] + prod[344][3447] + prod[345][3457] + prod[346][3467] + prod[347][3477] + prod[348][3487] + prod[349][3497] + prod[350][3507] + prod[351][3517] + prod[352][3527] + prod[353][3537] + prod[354][3547] + prod[355][3557] + prod[356][3567] + prod[357][3577] + prod[358][3587] + prod[359][3597] + prod[360][3607] + prod[361][3617] + prod[362][3627] + prod[363][3637] + prod[364][3647] + prod[365][3657] + prod[366][3667] + prod[367][3677] + prod[368][3687] + prod[369][3697] + prod[370][3707] + prod[371][3717] + prod[372][3727] + prod[373][3737] + prod[374][3747] + prod[375][3757] + prod[376][3767] + prod[377][3777] + prod[378][3787] + prod[379][3797] + prod[380][3807] + prod[381][3817] + prod[382][3827] + prod[383][3837] + prod[384][3847] + prod[385][3857] + prod[386][3867] + prod[387][3877] + prod[388][3887] + prod[389][3897] + prod[390][3907] + prod[391][3917] + prod[392][3927] + prod[393][3937] + prod[394][3947] + prod[395][3957] + prod[396][3967] + prod[397][3977] + prod[398][3987] + prod[399][3997] + prod[400][4007] + prod[401][4017] + prod[402][4027] + prod[403][4037] + prod[404][4047] + prod[405][4057] + prod[406][4067] + prod[407][4077] + prod[408][4087] + prod[409][4097] + prod[410][4107] + prod[411][4117] + prod[412][4127] + prod[413][4137] + prod[414][4147] + prod[415][4157] + prod[416][4167] + prod[417][4177] + prod[418][4187] + prod[419][4197] + prod[420][4207] + prod[421][4217] + prod[422][4227] + prod[423][4237] + prod[424][4247] + prod[425][4257] + prod[426][4267] + prod[427][4277] + prod[428][4287] + prod[429][4297] + prod[430][4307] + prod[431][4317] + prod[432][4327] + prod[433][4337] + prod[434][4347] + prod[435][4357] + prod[436][4367] + prod[437][4377] + prod[438][4387] + prod[439][4397] + prod[440][4407] + prod[441][4417] + prod[442][4427] + prod[443][4437] + prod[444][4447] + prod[445][4457] + prod[446][4467] + prod[447][4477] + prod[448][4487] + prod[449][4497] + prod[450][4507] + prod[451][4517] + prod[452][4527] + prod[453][4537] + prod[454][4547] + prod[455][4557] + prod[456][4567] + prod[457][4577] + prod[458][4587] + prod[459][4597] + prod[460][4607] + prod[461][4617] + prod[462][4627] + prod[463][4637] + prod[464][4647] + prod[465][4657] + prod[466][4667] + prod[467][4677] + prod[468][4687] + prod[469][4697] + prod[470][4707] + prod[471][4717] + prod[472][4727] + prod[473][4737] + prod[474][4747] + prod[475][4757] + prod[476][4767] + prod[477][4777] + prod[478][4787] + prod[479][4797] + prod[480][4807] + prod[481][4817] + prod[482][4827] + prod[483][4837] + prod[484][4847] + prod[485][4857] + prod[486][4867] + prod[487][4877] + prod[488][4887] + prod[489][4897] + prod[490][4907] + prod[491][4917] + prod[492][4927] + prod[493][4937] + prod[494][4947] + prod[495][4957] + prod[496][4967] + prod[497][4977] + prod[498][4987] + prod[499][4997] + prod[500][5007] + prod[501][5017] + prod[502][5027] + prod[503][5037] + prod[504][5047] + prod[505][5057] + prod[506][5067] + prod[507][5077] + prod[508][5087] + prod[509][5097] + prod[510][5107] + prod[511][5117] + prod[512][5127] + prod[513][5137] + prod[514][5147] + prod[515][5157] + prod[516][5167] + prod[517][5177] + prod[518][5187] + prod[519][5197] + prod[520][5207] + prod[521][5217] + prod[522][5227] + prod[523][5237] + prod[524][5247] + prod[525][5257] + prod[526][5267] + prod[527][5277] + prod[528][5287] + prod[529][5297] + prod[530][5307] + prod[531][5317] + prod[532][5327] + prod[533][5337] + prod[534][5347] + prod[535][5357] + prod[536][5367] + prod[537][5377] + prod[538][5387] + prod[539][5397] + prod[540][5407] + prod[541][5417] + prod[542][5427] + prod[543][5437] + prod[544][5447] + prod[545][5457] + prod[546][5467] + prod[547][5477] + prod[548][5487] + prod[549][5497] + prod[550][5507] + prod[551][5517] + prod[552][5527] + prod[553][5537] + prod[554][5547] + prod[555][5557] + prod[556][5567] + prod[557][5577] + prod[558][5587] + prod[559][5597] + prod[560][5607] + prod[561][5617] + prod[562][5627] + prod[563][5637] + prod[564][5647] + prod[565][5657] + prod[566][5667] + prod[567][5677] + prod[568][5687] + prod[569][5697] + prod[570][5707] + prod[571][5717] + prod[572][5727] + prod[573][5737] + prod[574][5747] + prod[575][5757] + prod[576][5767] + prod[577][5777] + prod[578][5787] + prod[579][5797] + prod[580][5807] + prod[581][5817] + prod[582][5827] + prod[583][5837] + prod[584][5847] + prod[585][5857] + prod[586][5867] + prod[587][5877] + prod[588][5887] + prod[589][5897] + prod[590][5907] + prod[591][5917] + prod[592][5927] + prod[593][5937] + prod[594][5947] + prod[595][5957] + prod[596][5967] + prod[597][5977] + prod[598][5987] + prod[599][5997] + prod[600][6007] + prod[601][6017] + prod[602][6027] + prod[603][6037] + prod[604][6047] + prod[605][6057] + prod[606][6067] + prod[607][6077] + prod[608][6087] + prod[609][6097] + prod[610][6107] + prod[611][6117] + prod[612][6127] + prod[613][6137] + prod[614][6147] + prod[615][6157] + prod[616][6167] + prod[617][6177] + prod[618][6187] + prod[619][6197] + prod[620][6207] + prod[621][6217] + prod[622][6227] + prod[623][6237] + prod[624][6247] + prod[625][6257] + prod[626][6267] + prod[627][6277] + prod[628][6287] + prod[629][6297] + prod[630][6307] + prod[631][6317] + prod[632][6327] + prod[633][6337] + prod[634][6347] + prod[635][6357] + prod[636][6367] + prod[637][6377] + prod[638][6387] + prod[639][6397] + prod[640][6407] + prod[641][6417] + prod[642][6427] + prod[643][6437] + prod[644][6447] + prod[645][6457] + prod[646][6467] + prod[647][6477] + prod[648][6487] + prod[649][6497] + prod[650][6507] + prod[651][6517] + prod[652][6527] + prod[653][6537] + prod[654][6547] + prod[655][6557] + prod[656][6567] + prod[657][6577] + prod[658][6587] + prod[659][6597] + prod[660][6607] + prod[661][6617] + prod[662][6627] + prod[663][6637] + prod[664][6647] + prod[665][6657] + prod[666][6667] + prod[667][6677] + prod[668][6687] + prod[669][6697] + prod[670][6707] + prod[671][6717] + prod[672][6727] + prod[673][6737] + prod[674][6747] + prod[675][6757] + prod[676][6767] + prod[677][6777] + prod[678][6787] + prod[679][6797] + prod[680][6807] + prod[681][6817] + prod[682][6827] + prod[683][6837] + prod[684][6847] + prod[685][6857] + prod[686][6867] + prod[687][6877] + prod[688][6887] + prod[689][6897] + prod[690][6907] + prod[691][6917] + prod[692][6927] + prod[693][6937] + prod[694][6947] + prod[695][6957] + prod[696][6967] + prod[697][6977] + prod[698][6987] + prod[699][6997] + prod[700][7007] + prod[701][7017] + prod[702][7027] + prod[703][7037] + prod[704][7047] + prod[705][7057] + prod[706][7067] + prod[707][7077] + prod[708][7087] + prod[709][7097] + prod[710][7107] + prod[711][7117] + prod[712][7127] + prod[713][7137] + prod[714][7147] + prod[715][7157] + prod[716][7167] + prod[717][7177] + prod[718][7187] + prod[719][7197] + prod[720][7207] + prod[721][7217] + prod[722][7227] + prod[723][7237] + prod[724][7247] + prod[725][7257] + prod[726][7267] + prod[727][7277] + prod[728][7287] + prod[729][7297] + prod[730][7307] + prod[731][7317] + prod[732][7327] + prod[733][7337] + prod[734][7347] + prod[735][7357] + prod[736][7367] + prod[737][7377] + prod[738][7387] + prod[739][7397] + prod[740][7407] + prod[741][7417] + prod[742][7427] + prod[743][7437] + prod[744][7447] + prod[745][7457] + prod[746][7467] + prod[747][7477] + prod[748][7487] + prod[749][7497] + prod[750][7507] + prod[751][7517] + prod[752][7527] + prod[753][7537] + prod[754][7547] + prod[755][7557] + prod[756][7567] + prod[757][7577] + prod[758][7587] + prod[759][7597] + prod[760][7607] + prod[761][7617] + prod[762][7627] + prod[763][7637] + prod[764][7647] + prod[765][7657] + prod[766][7667] + prod[767][7677] + prod[768][7687] + prod[769][7697] + prod[770][7707] + prod[771][7717] + prod[772][7727] + prod[773][7737] + prod[774][7747] + prod[775][7757] + prod[776][7767] + prod[777][7777] + prod[778][7787] + prod[779][7797] + prod[780][7807] + prod[781][7817] + prod[782][7827] + prod[783][7837];
mul_temp[8] = prod[0][8] + prod[1][18] + prod[2][28] + prod[3][38] + prod[4][48] + prod[5][58] + prod[6][68] + prod[7][78] + prod[8][88] + prod[9][98] + prod[10][108] + prod[11][118] + prod[12][128] + prod[13][138] + prod[14][148] + prod[15][158] + prod[16][168] + prod[17][178] + prod[18][188] + prod[19][198] + prod[20][208] + prod[21][218] + prod[22][228] + prod[23][238] + prod[24][248] + prod[25][258] + prod[26][268] + prod[27][278] + prod[28][288] + prod[29][298] + prod[30][308] + prod[31][318] + prod[32][328] + prod[33][338] + prod[34][348] + prod[35][358] + prod[36][368] + prod[37][378] + prod[38][388] + prod[39][398] + prod[40][408] + prod[41][418] + prod[42][428] + prod[43][438] + prod[44][448] + prod[45][458] + prod[46][468] + prod[47][478] + prod[48][488] + prod[49][498] + prod[50][508] + prod[51][518] + prod[52][528] + prod[53][538] + prod[54][548] + prod[55][558] + prod[56][568] + prod[57][578] + prod[58][588] + prod[59][598] + prod[60][608] + prod[61][618] + prod[62][628] + prod[63][638] + prod[64][648] + prod[65][658] + prod[66][668] + prod[67][678] + prod[68][688] + prod[69][698] + prod[70][708] + prod[71][718] + prod[72][728] + prod[73][738] + prod[74][748] + prod[75][758] + prod[76][768] + prod[77][778] + prod[78][788] + prod[79][798] + prod[80][808] + prod[81][818] + prod[82][828] + prod[83][838] + prod[84][848] + prod[85][858] + prod[86][868] + prod[87][878] + prod[88][888] + prod[89][898] + prod[90][908] + prod[91][918] + prod[92][928] + prod[93][938] + prod[94][948] + prod[95][958] + prod[96][968] + prod[97][978] + prod[98][988] + prod[99][998] + prod[100][1008] + prod[101][1018] + prod[102][1028] + prod[103][1038] + prod[104][1048] + prod[105][1058] + prod[106][1068] + prod[107][1078] + prod[108][1088] + prod[109][1098] + prod[110][1108] + prod[111][1118] + prod[112][1128] + prod[113][1138] + prod[114][1148] + prod[115][1158] + prod[116][1168] + prod[117][1178] + prod[118][1188] + prod[119][1198] + prod[120][1208] + prod[121][1218] + prod[122][1228] + prod[123][1238] + prod[124][1248] + prod[125][1258] + prod[126][1268] + prod[127][1278] + prod[128][1288] + prod[129][1298] + prod[130][1308] + prod[131][1318] + prod[132][1328] + prod[133][1338] + prod[134][1348] + prod[135][1358] + prod[136][1368] + prod[137][1378] + prod[138][1388] + prod[139][1398] + prod[140][1408] + prod[141][1418] + prod[142][1428] + prod[143][1438] + prod[144][1448] + prod[145][1458] + prod[146][1468] + prod[147][1478] + prod[148][1488] + prod[149][1498] + prod[150][1508] + prod[151][1518] + prod[152][1528] + prod[153][1538] + prod[154][1548] + prod[155][1558] + prod[156][1568] + prod[157][1578] + prod[158][1588] + prod[159][1598] + prod[160][1608] + prod[161][1618] + prod[162][1628] + prod[163][1638] + prod[164][1648] + prod[165][1658] + prod[166][1668] + prod[167][1678] + prod[168][1688] + prod[169][1698] + prod[170][1708] + prod[171][1718] + prod[172][1728] + prod[173][1738] + prod[174][1748] + prod[175][1758] + prod[176][1768] + prod[177][1778] + prod[178][1788] + prod[179][1798] + prod[180][1808] + prod[181][1818] + prod[182][1828] + prod[183][1838] + prod[184][1848] + prod[185][1858] + prod[186][1868] + prod[187][1878] + prod[188][1888] + prod[189][1898] + prod[190][1908] + prod[191][1918] + prod[192][1928] + prod[193][1938] + prod[194][1948] + prod[195][1958] + prod[196][1968] + prod[197][1978] + prod[198][1988] + prod[199][1998] + prod[200][2008] + prod[201][2018] + prod[202][2028] + prod[203][2038] + prod[204][2048] + prod[205][2058] + prod[206][2068] + prod[207][2078] + prod[208][2088] + prod[209][2098] + prod[210][2108] + prod[211][2118] + prod[212][2128] + prod[213][2138] + prod[214][2148] + prod[215][2158] + prod[216][2168] + prod[217][2178] + prod[218][2188] + prod[219][2198] + prod[220][2208] + prod[221][2218] + prod[222][2228] + prod[223][2238] + prod[224][2248] + prod[225][2258] + prod[226][2268] + prod[227][2278] + prod[228][2288] + prod[229][2298] + prod[230][2308] + prod[231][2318] + prod[232][2328] + prod[233][2338] + prod[234][2348] + prod[235][2358] + prod[236][2368] + prod[237][2378] + prod[238][2388] + prod[239][2398] + prod[240][2408] + prod[241][2418] + prod[242][2428] + prod[243][2438] + prod[244][2448] + prod[245][2458] + prod[246][2468] + prod[247][2478] + prod[248][2488] + prod[249][2498] + prod[250][2508] + prod[251][2518] + prod[252][2528] + prod[253][2538] + prod[254][2548] + prod[255][2558] + prod[256][2568] + prod[257][2578] + prod[258][2588] + prod[259][2598] + prod[260][2608] + prod[261][2618] + prod[262][2628] + prod[263][2638] + prod[264][2648] + prod[265][2658] + prod[266][2668] + prod[267][2678] + prod[268][2688] + prod[269][2698] + prod[270][2708] + prod[271][2718] + prod[272][2728] + prod[273][2738] + prod[274][2748] + prod[275][2758] + prod[276][2768] + prod[277][2778] + prod[278][2788] + prod[279][2798] + prod[280][2808] + prod[281][2818] + prod[282][2828] + prod[283][2838] + prod[284][2848] + prod[285][2858] + prod[286][2868] + prod[287][2878] + prod[288][2888] + prod[289][2898] + prod[290][2908] + prod[291][2918] + prod[292][2928] + prod[293][2938] + prod[294][2948] + prod[295][2958] + prod[296][2968] + prod[297][2978] + prod[298][2988] + prod[299][2998] + prod[300][3008] + prod[301][3018] + prod[302][3028] + prod[303][3038] + prod[304][3048] + prod[305][3058] + prod[306][3068] + prod[307][3078] + prod[308][3088] + prod[309][3098] + prod[310][3108] + prod[311][3118] + prod[312][3128] + prod[313][3138] + prod[314][3148] + prod[315][3158] + prod[316][3168] + prod[317][3178] + prod[318][3188] + prod[319][3198] + prod[320][3208] + prod[321][3218] + prod[322][3228] + prod[323][3238] + prod[324][3248] + prod[325][3258] + prod[326][3268] + prod[327][3278] + prod[328][3288] + prod[329][3298] + prod[330][3308] + prod[331][3318] + prod[332][3328] + prod[333][3338] + prod[334][3348] + prod[335][3358] + prod[336][3368] + prod[337][3378] + prod[338][3388] + prod[339][3398] + prod[340][3408] + prod[341][3418] + prod[342][3428] + prod[343][3438] + prod[344][3448] + prod[345][3458] + prod[346][3468] + prod[347][3478] + prod[348][3488] + prod[349][3498] + prod[350][3508] + prod[351][3518] + prod[352][3528] + prod[353][3538] + prod[354][3548] + prod[355][3558] + prod[356][3568] + prod[357][3578] + prod[358][3588] + prod[359][3598] + prod[360][3608] + prod[361][3618] + prod[362][3628] + prod[363][3638] + prod[364][3648] + prod[365][3658] + prod[366][3668] + prod[367][3678] + prod[368][3688] + prod[369][3698] + prod[370][3708] + prod[371][3718] + prod[372][3728] + prod[373][3738] + prod[374][3748] + prod[375][3758] + prod[376][3768] + prod[377][3778] + prod[378][3788] + prod[379][3798] + prod[380][3808] + prod[381][3818] + prod[382][3828] + prod[383][3838] + prod[384][3848] + prod[385][3858] + prod[386][3868] + prod[387][3878] + prod[388][3888] + prod[389][3898] + prod[390][3908] + prod[391][3918] + prod[392][3928] + prod[393][3938] + prod[394][3948] + prod[395][3958] + prod[396][3968] + prod[397][3978] + prod[398][3988] + prod[399][3998] + prod[400][4008] + prod[401][4018] + prod[402][4028] + prod[403][4038] + prod[404][4048] + prod[405][4058] + prod[406][4068] + prod[407][4078] + prod[408][4088] + prod[409][4098] + prod[410][4108] + prod[411][4118] + prod[412][4128] + prod[413][4138] + prod[414][4148] + prod[415][4158] + prod[416][4168] + prod[417][4178] + prod[418][4188] + prod[419][4198] + prod[420][4208] + prod[421][4218] + prod[422][4228] + prod[423][4238] + prod[424][4248] + prod[425][4258] + prod[426][4268] + prod[427][4278] + prod[428][4288] + prod[429][4298] + prod[430][4308] + prod[431][4318] + prod[432][4328] + prod[433][4338] + prod[434][4348] + prod[435][4358] + prod[436][4368] + prod[437][4378] + prod[438][4388] + prod[439][4398] + prod[440][4408] + prod[441][4418] + prod[442][4428] + prod[443][4438] + prod[444][4448] + prod[445][4458] + prod[446][4468] + prod[447][4478] + prod[448][4488] + prod[449][4498] + prod[450][4508] + prod[451][4518] + prod[452][4528] + prod[453][4538] + prod[454][4548] + prod[455][4558] + prod[456][4568] + prod[457][4578] + prod[458][4588] + prod[459][4598] + prod[460][4608] + prod[461][4618] + prod[462][4628] + prod[463][4638] + prod[464][4648] + prod[465][4658] + prod[466][4668] + prod[467][4678] + prod[468][4688] + prod[469][4698] + prod[470][4708] + prod[471][4718] + prod[472][4728] + prod[473][4738] + prod[474][4748] + prod[475][4758] + prod[476][4768] + prod[477][4778] + prod[478][4788] + prod[479][4798] + prod[480][4808] + prod[481][4818] + prod[482][4828] + prod[483][4838] + prod[484][4848] + prod[485][4858] + prod[486][4868] + prod[487][4878] + prod[488][4888] + prod[489][4898] + prod[490][4908] + prod[491][4918] + prod[492][4928] + prod[493][4938] + prod[494][4948] + prod[495][4958] + prod[496][4968] + prod[497][4978] + prod[498][4988] + prod[499][4998] + prod[500][5008] + prod[501][5018] + prod[502][5028] + prod[503][5038] + prod[504][5048] + prod[505][5058] + prod[506][5068] + prod[507][5078] + prod[508][5088] + prod[509][5098] + prod[510][5108] + prod[511][5118] + prod[512][5128] + prod[513][5138] + prod[514][5148] + prod[515][5158] + prod[516][5168] + prod[517][5178] + prod[518][5188] + prod[519][5198] + prod[520][5208] + prod[521][5218] + prod[522][5228] + prod[523][5238] + prod[524][5248] + prod[525][5258] + prod[526][5268] + prod[527][5278] + prod[528][5288] + prod[529][5298] + prod[530][5308] + prod[531][5318] + prod[532][5328] + prod[533][5338] + prod[534][5348] + prod[535][5358] + prod[536][5368] + prod[537][5378] + prod[538][5388] + prod[539][5398] + prod[540][5408] + prod[541][5418] + prod[542][5428] + prod[543][5438] + prod[544][5448] + prod[545][5458] + prod[546][5468] + prod[547][5478] + prod[548][5488] + prod[549][5498] + prod[550][5508] + prod[551][5518] + prod[552][5528] + prod[553][5538] + prod[554][5548] + prod[555][5558] + prod[556][5568] + prod[557][5578] + prod[558][5588] + prod[559][5598] + prod[560][5608] + prod[561][5618] + prod[562][5628] + prod[563][5638] + prod[564][5648] + prod[565][5658] + prod[566][5668] + prod[567][5678] + prod[568][5688] + prod[569][5698] + prod[570][5708] + prod[571][5718] + prod[572][5728] + prod[573][5738] + prod[574][5748] + prod[575][5758] + prod[576][5768] + prod[577][5778] + prod[578][5788] + prod[579][5798] + prod[580][5808] + prod[581][5818] + prod[582][5828] + prod[583][5838] + prod[584][5848] + prod[585][5858] + prod[586][5868] + prod[587][5878] + prod[588][5888] + prod[589][5898] + prod[590][5908] + prod[591][5918] + prod[592][5928] + prod[593][5938] + prod[594][5948] + prod[595][5958] + prod[596][5968] + prod[597][5978] + prod[598][5988] + prod[599][5998] + prod[600][6008] + prod[601][6018] + prod[602][6028] + prod[603][6038] + prod[604][6048] + prod[605][6058] + prod[606][6068] + prod[607][6078] + prod[608][6088] + prod[609][6098] + prod[610][6108] + prod[611][6118] + prod[612][6128] + prod[613][6138] + prod[614][6148] + prod[615][6158] + prod[616][6168] + prod[617][6178] + prod[618][6188] + prod[619][6198] + prod[620][6208] + prod[621][6218] + prod[622][6228] + prod[623][6238] + prod[624][6248] + prod[625][6258] + prod[626][6268] + prod[627][6278] + prod[628][6288] + prod[629][6298] + prod[630][6308] + prod[631][6318] + prod[632][6328] + prod[633][6338] + prod[634][6348] + prod[635][6358] + prod[636][6368] + prod[637][6378] + prod[638][6388] + prod[639][6398] + prod[640][6408] + prod[641][6418] + prod[642][6428] + prod[643][6438] + prod[644][6448] + prod[645][6458] + prod[646][6468] + prod[647][6478] + prod[648][6488] + prod[649][6498] + prod[650][6508] + prod[651][6518] + prod[652][6528] + prod[653][6538] + prod[654][6548] + prod[655][6558] + prod[656][6568] + prod[657][6578] + prod[658][6588] + prod[659][6598] + prod[660][6608] + prod[661][6618] + prod[662][6628] + prod[663][6638] + prod[664][6648] + prod[665][6658] + prod[666][6668] + prod[667][6678] + prod[668][6688] + prod[669][6698] + prod[670][6708] + prod[671][6718] + prod[672][6728] + prod[673][6738] + prod[674][6748] + prod[675][6758] + prod[676][6768] + prod[677][6778] + prod[678][6788] + prod[679][6798] + prod[680][6808] + prod[681][6818] + prod[682][6828] + prod[683][6838] + prod[684][6848] + prod[685][6858] + prod[686][6868] + prod[687][6878] + prod[688][6888] + prod[689][6898] + prod[690][6908] + prod[691][6918] + prod[692][6928] + prod[693][6938] + prod[694][6948] + prod[695][6958] + prod[696][6968] + prod[697][6978] + prod[698][6988] + prod[699][6998] + prod[700][7008] + prod[701][7018] + prod[702][7028] + prod[703][7038] + prod[704][7048] + prod[705][7058] + prod[706][7068] + prod[707][7078] + prod[708][7088] + prod[709][7098] + prod[710][7108] + prod[711][7118] + prod[712][7128] + prod[713][7138] + prod[714][7148] + prod[715][7158] + prod[716][7168] + prod[717][7178] + prod[718][7188] + prod[719][7198] + prod[720][7208] + prod[721][7218] + prod[722][7228] + prod[723][7238] + prod[724][7248] + prod[725][7258] + prod[726][7268] + prod[727][7278] + prod[728][7288] + prod[729][7298] + prod[730][7308] + prod[731][7318] + prod[732][7328] + prod[733][7338] + prod[734][7348] + prod[735][7358] + prod[736][7368] + prod[737][7378] + prod[738][7388] + prod[739][7398] + prod[740][7408] + prod[741][7418] + prod[742][7428] + prod[743][7438] + prod[744][7448] + prod[745][7458] + prod[746][7468] + prod[747][7478] + prod[748][7488] + prod[749][7498] + prod[750][7508] + prod[751][7518] + prod[752][7528] + prod[753][7538] + prod[754][7548] + prod[755][7558] + prod[756][7568] + prod[757][7578] + prod[758][7588] + prod[759][7598] + prod[760][7608] + prod[761][7618] + prod[762][7628] + prod[763][7638] + prod[764][7648] + prod[765][7658] + prod[766][7668] + prod[767][7678] + prod[768][7688] + prod[769][7698] + prod[770][7708] + prod[771][7718] + prod[772][7728] + prod[773][7738] + prod[774][7748] + prod[775][7758] + prod[776][7768] + prod[777][7778] + prod[778][7788] + prod[779][7798] + prod[780][7808] + prod[781][7818] + prod[782][7828] + prod[783][7838];
mul_temp[9] = prod[0][9] + prod[1][19] + prod[2][29] + prod[3][39] + prod[4][49] + prod[5][59] + prod[6][69] + prod[7][79] + prod[8][89] + prod[9][99] + prod[10][109] + prod[11][119] + prod[12][129] + prod[13][139] + prod[14][149] + prod[15][159] + prod[16][169] + prod[17][179] + prod[18][189] + prod[19][199] + prod[20][209] + prod[21][219] + prod[22][229] + prod[23][239] + prod[24][249] + prod[25][259] + prod[26][269] + prod[27][279] + prod[28][289] + prod[29][299] + prod[30][309] + prod[31][319] + prod[32][329] + prod[33][339] + prod[34][349] + prod[35][359] + prod[36][369] + prod[37][379] + prod[38][389] + prod[39][399] + prod[40][409] + prod[41][419] + prod[42][429] + prod[43][439] + prod[44][449] + prod[45][459] + prod[46][469] + prod[47][479] + prod[48][489] + prod[49][499] + prod[50][509] + prod[51][519] + prod[52][529] + prod[53][539] + prod[54][549] + prod[55][559] + prod[56][569] + prod[57][579] + prod[58][589] + prod[59][599] + prod[60][609] + prod[61][619] + prod[62][629] + prod[63][639] + prod[64][649] + prod[65][659] + prod[66][669] + prod[67][679] + prod[68][689] + prod[69][699] + prod[70][709] + prod[71][719] + prod[72][729] + prod[73][739] + prod[74][749] + prod[75][759] + prod[76][769] + prod[77][779] + prod[78][789] + prod[79][799] + prod[80][809] + prod[81][819] + prod[82][829] + prod[83][839] + prod[84][849] + prod[85][859] + prod[86][869] + prod[87][879] + prod[88][889] + prod[89][899] + prod[90][909] + prod[91][919] + prod[92][929] + prod[93][939] + prod[94][949] + prod[95][959] + prod[96][969] + prod[97][979] + prod[98][989] + prod[99][999] + prod[100][1009] + prod[101][1019] + prod[102][1029] + prod[103][1039] + prod[104][1049] + prod[105][1059] + prod[106][1069] + prod[107][1079] + prod[108][1089] + prod[109][1099] + prod[110][1109] + prod[111][1119] + prod[112][1129] + prod[113][1139] + prod[114][1149] + prod[115][1159] + prod[116][1169] + prod[117][1179] + prod[118][1189] + prod[119][1199] + prod[120][1209] + prod[121][1219] + prod[122][1229] + prod[123][1239] + prod[124][1249] + prod[125][1259] + prod[126][1269] + prod[127][1279] + prod[128][1289] + prod[129][1299] + prod[130][1309] + prod[131][1319] + prod[132][1329] + prod[133][1339] + prod[134][1349] + prod[135][1359] + prod[136][1369] + prod[137][1379] + prod[138][1389] + prod[139][1399] + prod[140][1409] + prod[141][1419] + prod[142][1429] + prod[143][1439] + prod[144][1449] + prod[145][1459] + prod[146][1469] + prod[147][1479] + prod[148][1489] + prod[149][1499] + prod[150][1509] + prod[151][1519] + prod[152][1529] + prod[153][1539] + prod[154][1549] + prod[155][1559] + prod[156][1569] + prod[157][1579] + prod[158][1589] + prod[159][1599] + prod[160][1609] + prod[161][1619] + prod[162][1629] + prod[163][1639] + prod[164][1649] + prod[165][1659] + prod[166][1669] + prod[167][1679] + prod[168][1689] + prod[169][1699] + prod[170][1709] + prod[171][1719] + prod[172][1729] + prod[173][1739] + prod[174][1749] + prod[175][1759] + prod[176][1769] + prod[177][1779] + prod[178][1789] + prod[179][1799] + prod[180][1809] + prod[181][1819] + prod[182][1829] + prod[183][1839] + prod[184][1849] + prod[185][1859] + prod[186][1869] + prod[187][1879] + prod[188][1889] + prod[189][1899] + prod[190][1909] + prod[191][1919] + prod[192][1929] + prod[193][1939] + prod[194][1949] + prod[195][1959] + prod[196][1969] + prod[197][1979] + prod[198][1989] + prod[199][1999] + prod[200][2009] + prod[201][2019] + prod[202][2029] + prod[203][2039] + prod[204][2049] + prod[205][2059] + prod[206][2069] + prod[207][2079] + prod[208][2089] + prod[209][2099] + prod[210][2109] + prod[211][2119] + prod[212][2129] + prod[213][2139] + prod[214][2149] + prod[215][2159] + prod[216][2169] + prod[217][2179] + prod[218][2189] + prod[219][2199] + prod[220][2209] + prod[221][2219] + prod[222][2229] + prod[223][2239] + prod[224][2249] + prod[225][2259] + prod[226][2269] + prod[227][2279] + prod[228][2289] + prod[229][2299] + prod[230][2309] + prod[231][2319] + prod[232][2329] + prod[233][2339] + prod[234][2349] + prod[235][2359] + prod[236][2369] + prod[237][2379] + prod[238][2389] + prod[239][2399] + prod[240][2409] + prod[241][2419] + prod[242][2429] + prod[243][2439] + prod[244][2449] + prod[245][2459] + prod[246][2469] + prod[247][2479] + prod[248][2489] + prod[249][2499] + prod[250][2509] + prod[251][2519] + prod[252][2529] + prod[253][2539] + prod[254][2549] + prod[255][2559] + prod[256][2569] + prod[257][2579] + prod[258][2589] + prod[259][2599] + prod[260][2609] + prod[261][2619] + prod[262][2629] + prod[263][2639] + prod[264][2649] + prod[265][2659] + prod[266][2669] + prod[267][2679] + prod[268][2689] + prod[269][2699] + prod[270][2709] + prod[271][2719] + prod[272][2729] + prod[273][2739] + prod[274][2749] + prod[275][2759] + prod[276][2769] + prod[277][2779] + prod[278][2789] + prod[279][2799] + prod[280][2809] + prod[281][2819] + prod[282][2829] + prod[283][2839] + prod[284][2849] + prod[285][2859] + prod[286][2869] + prod[287][2879] + prod[288][2889] + prod[289][2899] + prod[290][2909] + prod[291][2919] + prod[292][2929] + prod[293][2939] + prod[294][2949] + prod[295][2959] + prod[296][2969] + prod[297][2979] + prod[298][2989] + prod[299][2999] + prod[300][3009] + prod[301][3019] + prod[302][3029] + prod[303][3039] + prod[304][3049] + prod[305][3059] + prod[306][3069] + prod[307][3079] + prod[308][3089] + prod[309][3099] + prod[310][3109] + prod[311][3119] + prod[312][3129] + prod[313][3139] + prod[314][3149] + prod[315][3159] + prod[316][3169] + prod[317][3179] + prod[318][3189] + prod[319][3199] + prod[320][3209] + prod[321][3219] + prod[322][3229] + prod[323][3239] + prod[324][3249] + prod[325][3259] + prod[326][3269] + prod[327][3279] + prod[328][3289] + prod[329][3299] + prod[330][3309] + prod[331][3319] + prod[332][3329] + prod[333][3339] + prod[334][3349] + prod[335][3359] + prod[336][3369] + prod[337][3379] + prod[338][3389] + prod[339][3399] + prod[340][3409] + prod[341][3419] + prod[342][3429] + prod[343][3439] + prod[344][3449] + prod[345][3459] + prod[346][3469] + prod[347][3479] + prod[348][3489] + prod[349][3499] + prod[350][3509] + prod[351][3519] + prod[352][3529] + prod[353][3539] + prod[354][3549] + prod[355][3559] + prod[356][3569] + prod[357][3579] + prod[358][3589] + prod[359][3599] + prod[360][3609] + prod[361][3619] + prod[362][3629] + prod[363][3639] + prod[364][3649] + prod[365][3659] + prod[366][3669] + prod[367][3679] + prod[368][3689] + prod[369][3699] + prod[370][3709] + prod[371][3719] + prod[372][3729] + prod[373][3739] + prod[374][3749] + prod[375][3759] + prod[376][3769] + prod[377][3779] + prod[378][3789] + prod[379][3799] + prod[380][3809] + prod[381][3819] + prod[382][3829] + prod[383][3839] + prod[384][3849] + prod[385][3859] + prod[386][3869] + prod[387][3879] + prod[388][3889] + prod[389][3899] + prod[390][3909] + prod[391][3919] + prod[392][3929] + prod[393][3939] + prod[394][3949] + prod[395][3959] + prod[396][3969] + prod[397][3979] + prod[398][3989] + prod[399][3999] + prod[400][4009] + prod[401][4019] + prod[402][4029] + prod[403][4039] + prod[404][4049] + prod[405][4059] + prod[406][4069] + prod[407][4079] + prod[408][4089] + prod[409][4099] + prod[410][4109] + prod[411][4119] + prod[412][4129] + prod[413][4139] + prod[414][4149] + prod[415][4159] + prod[416][4169] + prod[417][4179] + prod[418][4189] + prod[419][4199] + prod[420][4209] + prod[421][4219] + prod[422][4229] + prod[423][4239] + prod[424][4249] + prod[425][4259] + prod[426][4269] + prod[427][4279] + prod[428][4289] + prod[429][4299] + prod[430][4309] + prod[431][4319] + prod[432][4329] + prod[433][4339] + prod[434][4349] + prod[435][4359] + prod[436][4369] + prod[437][4379] + prod[438][4389] + prod[439][4399] + prod[440][4409] + prod[441][4419] + prod[442][4429] + prod[443][4439] + prod[444][4449] + prod[445][4459] + prod[446][4469] + prod[447][4479] + prod[448][4489] + prod[449][4499] + prod[450][4509] + prod[451][4519] + prod[452][4529] + prod[453][4539] + prod[454][4549] + prod[455][4559] + prod[456][4569] + prod[457][4579] + prod[458][4589] + prod[459][4599] + prod[460][4609] + prod[461][4619] + prod[462][4629] + prod[463][4639] + prod[464][4649] + prod[465][4659] + prod[466][4669] + prod[467][4679] + prod[468][4689] + prod[469][4699] + prod[470][4709] + prod[471][4719] + prod[472][4729] + prod[473][4739] + prod[474][4749] + prod[475][4759] + prod[476][4769] + prod[477][4779] + prod[478][4789] + prod[479][4799] + prod[480][4809] + prod[481][4819] + prod[482][4829] + prod[483][4839] + prod[484][4849] + prod[485][4859] + prod[486][4869] + prod[487][4879] + prod[488][4889] + prod[489][4899] + prod[490][4909] + prod[491][4919] + prod[492][4929] + prod[493][4939] + prod[494][4949] + prod[495][4959] + prod[496][4969] + prod[497][4979] + prod[498][4989] + prod[499][4999] + prod[500][5009] + prod[501][5019] + prod[502][5029] + prod[503][5039] + prod[504][5049] + prod[505][5059] + prod[506][5069] + prod[507][5079] + prod[508][5089] + prod[509][5099] + prod[510][5109] + prod[511][5119] + prod[512][5129] + prod[513][5139] + prod[514][5149] + prod[515][5159] + prod[516][5169] + prod[517][5179] + prod[518][5189] + prod[519][5199] + prod[520][5209] + prod[521][5219] + prod[522][5229] + prod[523][5239] + prod[524][5249] + prod[525][5259] + prod[526][5269] + prod[527][5279] + prod[528][5289] + prod[529][5299] + prod[530][5309] + prod[531][5319] + prod[532][5329] + prod[533][5339] + prod[534][5349] + prod[535][5359] + prod[536][5369] + prod[537][5379] + prod[538][5389] + prod[539][5399] + prod[540][5409] + prod[541][5419] + prod[542][5429] + prod[543][5439] + prod[544][5449] + prod[545][5459] + prod[546][5469] + prod[547][5479] + prod[548][5489] + prod[549][5499] + prod[550][5509] + prod[551][5519] + prod[552][5529] + prod[553][5539] + prod[554][5549] + prod[555][5559] + prod[556][5569] + prod[557][5579] + prod[558][5589] + prod[559][5599] + prod[560][5609] + prod[561][5619] + prod[562][5629] + prod[563][5639] + prod[564][5649] + prod[565][5659] + prod[566][5669] + prod[567][5679] + prod[568][5689] + prod[569][5699] + prod[570][5709] + prod[571][5719] + prod[572][5729] + prod[573][5739] + prod[574][5749] + prod[575][5759] + prod[576][5769] + prod[577][5779] + prod[578][5789] + prod[579][5799] + prod[580][5809] + prod[581][5819] + prod[582][5829] + prod[583][5839] + prod[584][5849] + prod[585][5859] + prod[586][5869] + prod[587][5879] + prod[588][5889] + prod[589][5899] + prod[590][5909] + prod[591][5919] + prod[592][5929] + prod[593][5939] + prod[594][5949] + prod[595][5959] + prod[596][5969] + prod[597][5979] + prod[598][5989] + prod[599][5999] + prod[600][6009] + prod[601][6019] + prod[602][6029] + prod[603][6039] + prod[604][6049] + prod[605][6059] + prod[606][6069] + prod[607][6079] + prod[608][6089] + prod[609][6099] + prod[610][6109] + prod[611][6119] + prod[612][6129] + prod[613][6139] + prod[614][6149] + prod[615][6159] + prod[616][6169] + prod[617][6179] + prod[618][6189] + prod[619][6199] + prod[620][6209] + prod[621][6219] + prod[622][6229] + prod[623][6239] + prod[624][6249] + prod[625][6259] + prod[626][6269] + prod[627][6279] + prod[628][6289] + prod[629][6299] + prod[630][6309] + prod[631][6319] + prod[632][6329] + prod[633][6339] + prod[634][6349] + prod[635][6359] + prod[636][6369] + prod[637][6379] + prod[638][6389] + prod[639][6399] + prod[640][6409] + prod[641][6419] + prod[642][6429] + prod[643][6439] + prod[644][6449] + prod[645][6459] + prod[646][6469] + prod[647][6479] + prod[648][6489] + prod[649][6499] + prod[650][6509] + prod[651][6519] + prod[652][6529] + prod[653][6539] + prod[654][6549] + prod[655][6559] + prod[656][6569] + prod[657][6579] + prod[658][6589] + prod[659][6599] + prod[660][6609] + prod[661][6619] + prod[662][6629] + prod[663][6639] + prod[664][6649] + prod[665][6659] + prod[666][6669] + prod[667][6679] + prod[668][6689] + prod[669][6699] + prod[670][6709] + prod[671][6719] + prod[672][6729] + prod[673][6739] + prod[674][6749] + prod[675][6759] + prod[676][6769] + prod[677][6779] + prod[678][6789] + prod[679][6799] + prod[680][6809] + prod[681][6819] + prod[682][6829] + prod[683][6839] + prod[684][6849] + prod[685][6859] + prod[686][6869] + prod[687][6879] + prod[688][6889] + prod[689][6899] + prod[690][6909] + prod[691][6919] + prod[692][6929] + prod[693][6939] + prod[694][6949] + prod[695][6959] + prod[696][6969] + prod[697][6979] + prod[698][6989] + prod[699][6999] + prod[700][7009] + prod[701][7019] + prod[702][7029] + prod[703][7039] + prod[704][7049] + prod[705][7059] + prod[706][7069] + prod[707][7079] + prod[708][7089] + prod[709][7099] + prod[710][7109] + prod[711][7119] + prod[712][7129] + prod[713][7139] + prod[714][7149] + prod[715][7159] + prod[716][7169] + prod[717][7179] + prod[718][7189] + prod[719][7199] + prod[720][7209] + prod[721][7219] + prod[722][7229] + prod[723][7239] + prod[724][7249] + prod[725][7259] + prod[726][7269] + prod[727][7279] + prod[728][7289] + prod[729][7299] + prod[730][7309] + prod[731][7319] + prod[732][7329] + prod[733][7339] + prod[734][7349] + prod[735][7359] + prod[736][7369] + prod[737][7379] + prod[738][7389] + prod[739][7399] + prod[740][7409] + prod[741][7419] + prod[742][7429] + prod[743][7439] + prod[744][7449] + prod[745][7459] + prod[746][7469] + prod[747][7479] + prod[748][7489] + prod[749][7499] + prod[750][7509] + prod[751][7519] + prod[752][7529] + prod[753][7539] + prod[754][7549] + prod[755][7559] + prod[756][7569] + prod[757][7579] + prod[758][7589] + prod[759][7599] + prod[760][7609] + prod[761][7619] + prod[762][7629] + prod[763][7639] + prod[764][7649] + prod[765][7659] + prod[766][7669] + prod[767][7679] + prod[768][7689] + prod[769][7699] + prod[770][7709] + prod[771][7719] + prod[772][7729] + prod[773][7739] + prod[774][7749] + prod[775][7759] + prod[776][7769] + prod[777][7779] + prod[778][7789] + prod[779][7799] + prod[780][7809] + prod[781][7819] + prod[782][7829] + prod[783][7839];
        end
    end
    
    always_comb begin
        mult <= mul_temp;
    end

endmodule
