////////////////////////////////////////////////////////////////////////////
// Author       : Jeneel / Prajyot
// Coursework   : ECE 751
// Module       : TLUT test-bench
// Description  : Test bench for TLUT with adder trees
////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns
`include "simd_cell.sv"
`include "DEF.sv"

module t_lut_tb ();

    logic   clk;
    logic   rst_n;
    logic   enable;
    logic   [`DIM_ROW1*`DIM_COL1-1:0][`INPUT_WIDTH-1:0]input_bin;
    logic   [`DIM_ROW2*`DIM_COL2-1:0][`WEIGHT_WIDTH-1:0]weight_bin;
    logic   [`DIM_ROW1*`DIM_COL2-1:0][`ACC_WIDTH-1:0]product;
    integer i=0;
    

    simd_cell t_lut
    (
        .clk(clk),    // Clock
        .rst_n(rst_n),  // Asynchronous reset active low
        .enable(enable),
        .input_bin(input_bin), // input in binary
        .weight_bin(weight_bin), // weight in binary
        .accumulated_mult(product)
    );

    always #5 clk = ~clk;

    initial
    begin
        clk = 1;
        rst_n = 0;
	    enable = 0;
	    input_bin  = {8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd84,8'd185,8'd159,8'd151,8'd60,8'd36,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd222,8'd254,8'd254,8'd254,8'd254,8'd241,8'd198,8'd198,8'd198,8'd198,8'd198,8'd198,8'd198,8'd198,8'd170,8'd52,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd67,8'd114,8'd72,8'd114,8'd163,8'd227,8'd254,8'd225,8'd254,8'd254,8'd254,8'd250,8'd229,8'd254,8'd254,8'd140,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd17,8'd66,8'd14,8'd67,8'd67,8'd67,8'd59,8'd21,8'd236,8'd254,8'd106,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd83,8'd253,8'd209,8'd18,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd22,8'd233,8'd255,8'd83,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd129,8'd254,8'd238,8'd44,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd59,8'd249,8'd254,8'd62,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd133,8'd254,8'd187,8'd5,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd9,8'd205,8'd248,8'd58,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd126,8'd254,8'd182,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd75,8'd251,8'd240,8'd57,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd19,8'd221,8'd254,8'd166,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd3,8'd203,8'd254,8'd219,8'd35,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd38,8'd254,8'd254,8'd77,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd224,8'd254,8'd115,8'd1,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd133,8'd254,8'd254,8'd52,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd61,8'd242,8'd254,8'd254,8'd52,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd121,8'd254,8'd254,8'd219,8'd40,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd121,8'd254,8'd207,8'd18,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0};
	    weight_bin = {8'd2,-8'd2,-8'd1,8'd2,-8'd4,8'd3,-8'd1,8'd2,8'd1,-8'd1,8'd1,8'd0,8'd2,-8'd2,8'd0,8'd0,8'd1,8'd0,8'd4,8'd1,-8'd2,-8'd3,-8'd1,-8'd2,-8'd1,8'd0,8'd3,8'd2,-8'd4,8'd3,8'd1,8'd4,8'd3,-8'd4,-8'd4,-8'd2,8'd4,-8'd1,8'd2,-8'd2,8'd5,-8'd2,8'd3,8'd0,-8'd3,8'd2,-8'd3,8'd1,-8'd2,-8'd1,-8'd4,-8'd2,8'd2,-8'd1,8'd5,8'd4,8'd0,-8'd3,8'd3,8'd1,-8'd3,8'd3,8'd3,8'd4,-8'd3,-8'd2,-8'd1,-8'd1,-8'd6,-8'd6,-8'd2,-8'd7,-8'd5,-8'd6,-8'd4,-8'd3,-8'd1,8'd1,-8'd5,8'd2,-8'd3,-8'd3,8'd0,-8'd1,8'd3,-8'd3,-8'd4,8'd3,-8'd1,8'd2,8'd1,-8'd4,-8'd1,-8'd4,-8'd11,-8'd11,-8'd8,-8'd9,-8'd12,-8'd14,-8'd10,-8'd16,-8'd16,-8'd16,-8'd18,-8'd16,-8'd4,-8'd3,8'd3,8'd1,8'd1,8'd3,8'd4,-8'd3,8'd1,8'd3,8'd3,8'd1,-8'd6,-8'd7,-8'd9,-8'd9,-8'd8,-8'd15,-8'd10,-8'd9,-8'd8,-8'd8,-8'd9,-8'd6,-8'd17,-8'd13,-8'd4,-8'd7,-8'd4,-8'd2,-8'd1,8'd0,-8'd3,-8'd4,-8'd2,-8'd1,-8'd3,8'd2,8'd0,-8'd4,-8'd5,-8'd6,-8'd10,-8'd13,-8'd14,-8'd3,8'd1,8'd17,8'd17,8'd22,8'd23,8'd27,8'd24,8'd10,-8'd2,8'd1,-8'd5,-8'd6,-8'd14,-8'd5,-8'd3,-8'd1,-8'd4,-8'd2,-8'd1,8'd2,-8'd1,-8'd3,-8'd3,-8'd8,-8'd14,-8'd17,-8'd11,8'd0,8'd4,8'd13,8'd13,8'd25,8'd27,8'd37,8'd23,8'd21,8'd20,8'd16,8'd12,-8'd10,-8'd21,-8'd12,-8'd2,-8'd4,8'd2,8'd3,8'd4,-8'd4,-8'd3,-8'd10,-8'd7,-8'd16,-8'd19,-8'd11,-8'd5,8'd2,8'd11,8'd11,8'd11,8'd20,8'd23,8'd39,8'd37,8'd26,8'd19,8'd10,8'd12,8'd10,-8'd20,-8'd14,-8'd10,-8'd3,8'd2,-8'd3,-8'd1,8'd2,-8'd5,-8'd7,-8'd13,-8'd20,-8'd13,-8'd12,-8'd1,8'd3,-8'd2,8'd2,8'd8,8'd12,8'd33,8'd36,8'd32,8'd15,8'd6,8'd6,8'd11,8'd18,-8'd12,-8'd17,-8'd1,-8'd2,8'd0,8'd2,8'd0,-8'd5,-8'd6,-8'd8,-8'd13,-8'd11,-8'd8,-8'd5,-8'd4,-8'd4,-8'd2,-8'd1,8'd7,8'd3,8'd21,8'd26,8'd37,8'd25,8'd7,8'd5,8'd14,8'd31,8'd0,-8'd16,-8'd6,8'd0,-8'd1,8'd1,8'd3,-8'd1,-8'd10,-8'd11,-8'd13,-8'd2,-8'd9,-8'd10,-8'd10,-8'd4,8'd3,-8'd3,-8'd18,-8'd30,-8'd30,8'd2,8'd24,8'd27,8'd25,8'd18,8'd29,8'd47,8'd22,-8'd7,-8'd5,8'd4,8'd1,8'd4,-8'd2,-8'd5,-8'd17,-8'd7,8'd4,-8'd4,-8'd4,-8'd6,-8'd1,8'd3,-8'd2,-8'd21,-8'd56,-8'd81,-8'd77,-8'd46,-8'd8,8'd17,8'd22,8'd33,8'd44,8'd55,8'd34,-8'd4,8'd0,-8'd1,-8'd3,-8'd3,8'd1,-8'd2,-8'd14,-8'd2,8'd6,8'd10,-8'd4,-8'd8,8'd3,8'd5,-8'd2,-8'd41,-8'd87,-8'd109,-8'd108,-8'd71,-8'd28,-8'd9,8'd5,8'd24,8'd50,8'd55,8'd30,-8'd4,8'd3,-8'd1,8'd2,8'd0,-8'd5,-8'd5,-8'd5,8'd6,8'd11,8'd12,8'd3,8'd0,8'd19,8'd9,-8'd13,-8'd61,-8'd97,-8'd110,-8'd106,-8'd74,-8'd37,-8'd35,-8'd21,8'd14,8'd44,8'd55,8'd32,-8'd1,8'd1,8'd4,8'd1,-8'd2,8'd4,-8'd4,-8'd2,8'd19,8'd29,8'd23,8'd9,8'd18,8'd24,8'd4,-8'd27,-8'd77,-8'd104,-8'd114,-8'd96,-8'd61,-8'd35,-8'd21,-8'd8,8'd8,8'd32,8'd49,8'd24,8'd4,-8'd3,-8'd2,-8'd4,8'd4,8'd1,-8'd2,-8'd1,8'd28,8'd25,8'd24,8'd21,8'd25,8'd29,-8'd14,-8'd56,-8'd98,-8'd112,-8'd116,-8'd84,-8'd52,-8'd15,-8'd7,-8'd5,8'd13,8'd23,8'd41,8'd21,8'd2,-8'd3,8'd3,-8'd2,-8'd4,8'd1,-8'd4,8'd4,8'd28,8'd39,8'd29,8'd17,8'd21,8'd23,-8'd29,-8'd82,-8'd121,-8'd113,-8'd98,-8'd68,-8'd25,-8'd4,-8'd1,8'd4,8'd13,8'd22,8'd21,8'd14,8'd3,8'd3,8'd4,-8'd4,8'd2,8'd1,-8'd11,-8'd1,8'd24,8'd34,8'd25,8'd23,8'd28,8'd18,-8'd22,-8'd88,-8'd110,-8'd105,-8'd79,-8'd29,-8'd3,8'd10,8'd8,8'd14,8'd10,8'd13,8'd13,8'd2,-8'd5,-8'd4,-8'd2,-8'd1,-8'd3,-8'd2,-8'd15,-8'd2,8'd17,8'd24,8'd18,8'd13,8'd36,8'd44,-8'd12,-8'd65,-8'd83,-8'd72,-8'd35,-8'd12,8'd5,8'd8,8'd1,-8'd1,8'd3,8'd10,8'd5,8'd0,-8'd4,8'd1,8'd1,8'd2,8'd1,-8'd1,-8'd12,-8'd3,8'd10,8'd18,8'd18,8'd17,8'd29,8'd46,8'd20,-8'd15,-8'd27,-8'd29,-8'd13,-8'd6,-8'd1,-8'd9,-8'd11,-8'd1,8'd1,-8'd1,-8'd2,8'd3,-8'd3,-8'd3,-8'd3,-8'd2,-8'd1,-8'd2,-8'd11,-8'd5,8'd7,8'd14,8'd11,8'd15,8'd28,8'd51,8'd36,8'd10,-8'd7,-8'd12,-8'd9,-8'd9,-8'd10,-8'd14,-8'd17,-8'd4,8'd1,-8'd5,-8'd1,-8'd2,-8'd4,-8'd2,8'd3,8'd2,8'd4,-8'd1,-8'd2,-8'd5,8'd6,8'd13,8'd20,8'd13,8'd21,8'd36,8'd46,8'd24,8'd6,8'd1,-8'd6,-8'd12,-8'd19,-8'd14,-8'd11,-8'd10,-8'd6,-8'd7,-8'd6,-8'd3,8'd1,8'd1,8'd3,8'd2,8'd2,8'd4,-8'd1,-8'd6,-8'd1,8'd13,8'd17,8'd23,8'd26,8'd23,8'd38,8'd31,8'd32,8'd18,8'd7,8'd1,-8'd9,-8'd16,-8'd12,-8'd12,-8'd13,-8'd12,-8'd6,-8'd1,-8'd1,8'd4,8'd4,8'd3,8'd2,-8'd4,8'd3,-8'd8,-8'd3,-8'd3,8'd8,8'd14,8'd24,8'd28,8'd35,8'd34,8'd31,8'd15,8'd8,-8'd5,-8'd5,-8'd18,-8'd24,-8'd16,-8'd13,-8'd1,-8'd4,-8'd4,-8'd3,8'd2,-8'd1,-8'd4,8'd1,8'd0,8'd2,-8'd3,-8'd5,-8'd1,-8'd12,-8'd6,-8'd6,-8'd8,-8'd6,8'd2,-8'd3,-8'd4,-8'd12,-8'd17,-8'd25,-8'd18,-8'd18,-8'd16,-8'd10,-8'd6,-8'd5,8'd2,-8'd2,8'd3,8'd3,-8'd3,-8'd3,-8'd2,8'd3,8'd0,-8'd3,-8'd2,-8'd5,-8'd11,-8'd24,-8'd25,-8'd26,-8'd26,-8'd31,-8'd30,-8'd24,-8'd23,-8'd18,-8'd17,-8'd13,-8'd3,-8'd1,8'd0,-8'd5,8'd2,8'd3,8'd1,-8'd2,8'd0,-8'd2,8'd4,8'd4,-8'd1,-8'd4,8'd1,8'd0,-8'd2,-8'd11,-8'd6,-8'd8,-8'd10,-8'd11,-8'd8,-8'd7,-8'd11,-8'd3,-8'd1,8'd1,8'd1,-8'd2,8'd2,8'd3,8'd2,-8'd3,-8'd2,8'd4,8'd3,8'd3,-8'd2,-8'd1,-8'd3,-8'd3,8'd3,-8'd4,-8'd1,8'd1,-8'd3,8'd1,-8'd2,8'd0,-8'd6,-8'd1,-8'd6,8'd2,8'd3,-8'd2,8'd0,-8'd3,-8'd3,-8'd2,-8'd2,8'd1,-8'd1,8'd0};
        
        #300;
        
//        if(product != {13'd30,13'd36,13'd42,13'd66,13'd81,13'd96,13'd90,13'd111,13'd132}) begin   
//            $display("test 1 SUCCESS");
//        end else begin
//            $display("test 2 FAILED");
//        end

	    //input_bin = {4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4};
	    //weight_bin = {4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1};
        //#30;
        //if(product == {13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12}) begin 
        //    $display("test 2 SUCCESS");
        //end else begin
        //    $display("test 2 FAILED");
        //end

        //#30;
	    @(negedge clk);
        rst_n = 1;
	   
	    #5;
	    @(negedge clk);
	    enable = 1;
	    @(posedge clk);
	
        for (i=0; i<50; i=i+1)
   		@(posedge clk) ; 
	
        $finish;
    end
endmodule
