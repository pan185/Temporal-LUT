////////////////////////////////////////////////////////////////////////////
// Author       : Jeneel / Prajyot
// Coursework   : ECE 751
// Module       : TLUT test-bench
// Description  : Test bench for TLUT with adder trees
////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns
`include "simd_cell.sv"
`include "DEF.sv"

module t_lut_tb ();

    logic   clk;
    logic   rst_n;
    logic   enable;
    logic   [`DIM_ROW1*`DIM_COL1-1:0][`INPUT_WIDTH-1:0]input_bin;
    logic   [`DIM_ROW2*`DIM_COL2-1:0][`WEIGHT_WIDTH-1:0]weight_bin;
    logic   [`DIM_ROW1*`DIM_COL2-1:0][`ACC_WIDTH-1:0]product;
    logic [`INPUT_WIDTH-1:0] count;
    logic finish;
    //integer i=0;
    integer write_data;
    

    simd_cell t_lut
    (
        .clk(clk),    // Clock
        .rst_n(rst_n),  // Asynchronous reset active low
        .enable(enable),
        .input_bin(input_bin), // input in binary
        .weight_bin(weight_bin), // weight in binary
        .accumulated_mult(product),
	.cntOut(count),
	.finish(finish)
    );

    always #1 clk = ~clk;

    initial
    begin
        clk    = 1;
        rst_n  = 0;
        enable = 0;
        
	//prajyotg: Adding parameters to write product into a file
        write_data = $fopen("write_out.txt");

	    //TODO :: read the txt file automatically
	    // Input = 7
	    //input_bin  = {8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd3,8'd18,8'd18,8'd18,8'd126,8'd136,8'd175,8'd26,8'd166,8'd255,8'd247,8'd127,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd30,8'd36,8'd94,8'd154,8'd170,8'd253,8'd253,8'd253,8'd253,8'd253,8'd225,8'd172,8'd253,8'd242,8'd195,8'd64,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd49,8'd238,8'd253,8'd253,8'd253,8'd253,8'd253,8'd253,8'd253,8'd253,8'd251,8'd93,8'd82,8'd82,8'd56,8'd39,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd18,8'd219,8'd253,8'd253,8'd253,8'd253,8'd253,8'd198,8'd182,8'd247,8'd241,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd80,8'd156,8'd107,8'd253,8'd253,8'd205,8'd11,8'd0,8'd43,8'd154,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd14,8'd1,8'd154,8'd253,8'd90,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd139,8'd253,8'd190,8'd2,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd190,8'd253,8'd70,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd35,8'd241,8'd225,8'd160,8'd108,8'd1,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd81,8'd240,8'd253,8'd253,8'd119,8'd25,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd45,8'd186,8'd253,8'd253,8'd150,8'd27,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd16,8'd93,8'd252,8'd253,8'd187,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd249,8'd253,8'd249,8'd64,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd46,8'd130,8'd183,8'd253,8'd253,8'd207,8'd2,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd39,8'd148,8'd229,8'd253,8'd253,8'd253,8'd250,8'd182,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd24,8'd114,8'd221,8'd253,8'd253,8'd253,8'd253,8'd201,8'd78,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd23,8'd66,8'd213,8'd253,8'd253,8'd253,8'd253,8'd198,8'd81,8'd2,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd18,8'd171,8'd219,8'd253,8'd253,8'd253,8'd253,8'd195,8'd80,8'd9,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd55,8'd172,8'd226,8'd253,8'd253,8'd253,8'd253,8'd244,8'd133,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd136,8'd253,8'd253,8'd253,8'd212,8'd135,8'd132,8'd16,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0};
	    input_bin  = {4'd3, 4'd3, 4'd3, 4'd3};
	    weight_bin = {-4'd2,-4'd2,-4'd2, -4'd2};
	    /**************************************************************************
	    * Adding in values of different weights:
	    * Please uncomment out single value for weight and run the simulation.
	    * ************************************************************************/
	    // 0
            // weight_bin={9'd2,-9'd2,-9'd1,9'd2,-9'd4,9'd3,-9'd1,9'd2,9'd1,-9'd1,9'd1,9'd0,9'd2,-9'd2,9'd0,9'd0,9'd1,9'd0,9'd4,9'd1,-9'd2,-9'd3,-9'd1,-9'd2,-9'd1,9'd0,9'd3,9'd2,-9'd4,9'd3,9'd1,9'd4,9'd3,-9'd4,-9'd4,-9'd2,9'd4,-9'd1,9'd2,-9'd2,9'd5,-9'd2,9'd3,9'd0,-9'd3,9'd2,-9'd3,9'd1,-9'd2,-9'd1,-9'd4,-9'd2,9'd2,-9'd1,9'd5,9'd4,9'd0,-9'd3,9'd3,9'd1,-9'd3,9'd3,9'd3,9'd4,-9'd3,-9'd2,-9'd1,-9'd1,-9'd6,-9'd6,-9'd2,-9'd7,-9'd5,-9'd6,-9'd4,-9'd3,-9'd1,9'd1,-9'd5,9'd2,-9'd3,-9'd3,9'd0,-9'd1,9'd3,-9'd3,-9'd4,9'd3,-9'd1,9'd2,9'd1,-9'd4,-9'd1,-9'd4,-9'd11,-9'd11,-9'd8,-9'd9,-9'd12,-9'd14,-9'd10,-9'd16,-9'd16,-9'd16,-9'd18,-9'd16,-9'd4,-9'd3,9'd3,9'd1,9'd1,9'd3,9'd4,-9'd3,9'd1,9'd3,9'd3,9'd1,-9'd6,-9'd7,-9'd9,-9'd9,-9'd8,-9'd15,-9'd10,-9'd9,-9'd8,-9'd8,-9'd9,-9'd6,-9'd17,-9'd13,-9'd4,-9'd7,-9'd4,-9'd2,-9'd1,9'd0,-9'd3,-9'd4,-9'd2,-9'd1,-9'd3,9'd2,9'd0,-9'd4,-9'd5,-9'd6,-9'd10,-9'd13,-9'd14,-9'd3,9'd1,9'd17,9'd17,9'd22,9'd23,9'd27,9'd24,9'd10,-9'd2,9'd1,-9'd5,-9'd6,-9'd14,-9'd5,-9'd3,-9'd1,-9'd4,-9'd2,-9'd1,9'd2,-9'd1,-9'd3,-9'd3,-9'd8,-9'd14,-9'd17,-9'd11,9'd0,9'd4,9'd13,9'd13,9'd25,9'd27,9'd37,9'd23,9'd21,9'd20,9'd16,9'd12,-9'd10,-9'd21,-9'd12,-9'd2,-9'd4,9'd2,9'd3,9'd4,-9'd4,-9'd3,-9'd10,-9'd7,-9'd16,-9'd19,-9'd11,-9'd5,9'd2,9'd11,9'd11,9'd11,9'd20,9'd23,9'd39,9'd37,9'd26,9'd19,9'd10,9'd12,9'd10,-9'd20,-9'd14,-9'd10,-9'd3,9'd2,-9'd3,-9'd1,9'd2,-9'd5,-9'd7,-9'd13,-9'd20,-9'd13,-9'd12,-9'd1,9'd3,-9'd2,9'd2,9'd8,9'd12,9'd33,9'd36,9'd32,9'd15,9'd6,9'd6,9'd11,9'd18,-9'd12,-9'd17,-9'd1,-9'd2,9'd0,9'd2,9'd0,-9'd5,-9'd6,-9'd8,-9'd13,-9'd11,-9'd8,-9'd5,-9'd4,-9'd4,-9'd2,-9'd1,9'd7,9'd3,9'd21,9'd26,9'd37,9'd25,9'd7,9'd5,9'd14,9'd31,9'd0,-9'd16,-9'd6,9'd0,-9'd1,9'd1,9'd3,-9'd1,-9'd10,-9'd11,-9'd13,-9'd2,-9'd9,-9'd10,-9'd10,-9'd4,9'd3,-9'd3,-9'd18,-9'd30,-9'd30,9'd2,9'd24,9'd27,9'd25,9'd18,9'd29,9'd47,9'd22,-9'd7,-9'd5,9'd4,9'd1,9'd4,-9'd2,-9'd5,-9'd17,-9'd7,9'd4,-9'd4,-9'd4,-9'd6,-9'd1,9'd3,-9'd2,-9'd21,-9'd56,-9'd81,-9'd77,-9'd46,-9'd8,9'd17,9'd22,9'd33,9'd44,9'd55,9'd34,-9'd4,9'd0,-9'd1,-9'd3,-9'd3,9'd1,-9'd2,-9'd14,-9'd2,9'd6,9'd10,-9'd4,-9'd8,9'd3,9'd5,-9'd2,-9'd41,-9'd87,-9'd109,-9'd108,-9'd71,-9'd28,-9'd9,9'd5,9'd24,9'd50,9'd55,9'd30,-9'd4,9'd3,-9'd1,9'd2,9'd0,-9'd5,-9'd5,-9'd5,9'd6,9'd11,9'd12,9'd3,9'd0,9'd19,9'd9,-9'd13,-9'd61,-9'd97,-9'd110,-9'd106,-9'd74,-9'd37,-9'd35,-9'd21,9'd14,9'd44,9'd55,9'd32,-9'd1,9'd1,9'd4,9'd1,-9'd2,9'd4,-9'd4,-9'd2,9'd19,9'd29,9'd23,9'd9,9'd18,9'd24,9'd4,-9'd27,-9'd77,-9'd104,-9'd114,-9'd96,-9'd61,-9'd35,-9'd21,-9'd8,9'd8,9'd32,9'd49,9'd24,9'd4,-9'd3,-9'd2,-9'd4,9'd4,9'd1,-9'd2,-9'd1,9'd28,9'd25,9'd24,9'd21,9'd25,9'd29,-9'd14,-9'd56,-9'd98,-9'd112,-9'd116,-9'd84,-9'd52,-9'd15,-9'd7,-9'd5,9'd13,9'd23,9'd41,9'd21,9'd2,-9'd3,9'd3,-9'd2,-9'd4,9'd1,-9'd4,9'd4,9'd28,9'd39,9'd29,9'd17,9'd21,9'd23,-9'd29,-9'd82,-9'd121,-9'd113,-9'd98,-9'd68,-9'd25,-9'd4,-9'd1,9'd4,9'd13,9'd22,9'd21,9'd14,9'd3,9'd3,9'd4,-9'd4,9'd2,9'd1,-9'd11,-9'd1,9'd24,9'd34,9'd25,9'd23,9'd28,9'd18,-9'd22,-9'd88,-9'd110,-9'd105,-9'd79,-9'd29,-9'd3,9'd10,9'd8,9'd14,9'd10,9'd13,9'd13,9'd2,-9'd5,-9'd4,-9'd2,-9'd1,-9'd3,-9'd2,-9'd15,-9'd2,9'd17,9'd24,9'd18,9'd13,9'd36,9'd44,-9'd12,-9'd65,-9'd83,-9'd72,-9'd35,-9'd12,9'd5,9'd8,9'd1,-9'd1,9'd3,9'd10,9'd5,9'd0,-9'd4,9'd1,9'd1,9'd2,9'd1,-9'd1,-9'd12,-9'd3,9'd10,9'd18,9'd18,9'd17,9'd29,9'd46,9'd20,-9'd15,-9'd27,-9'd29,-9'd13,-9'd6,-9'd1,-9'd9,-9'd11,-9'd1,9'd1,-9'd1,-9'd2,9'd3,-9'd3,-9'd3,-9'd3,-9'd2,-9'd1,-9'd2,-9'd11,-9'd5,9'd7,9'd14,9'd11,9'd15,9'd28,9'd51,9'd36,9'd10,-9'd7,-9'd12,-9'd9,-9'd9,-9'd10,-9'd14,-9'd17,-9'd4,9'd1,-9'd5,-9'd1,-9'd2,-9'd4,-9'd2,9'd3,9'd2,9'd4,-9'd1,-9'd2,-9'd5,9'd6,9'd13,9'd20,9'd13,9'd21,9'd36,9'd46,9'd24,9'd6,9'd1,-9'd6,-9'd12,-9'd19,-9'd14,-9'd11,-9'd10,-9'd6,-9'd7,-9'd6,-9'd3,9'd1,9'd1,9'd3,9'd2,9'd2,9'd4,-9'd1,-9'd6,-9'd1,9'd13,9'd17,9'd23,9'd26,9'd23,9'd38,9'd31,9'd32,9'd18,9'd7,9'd1,-9'd9,-9'd16,-9'd12,-9'd12,-9'd13,-9'd12,-9'd6,-9'd1,-9'd1,9'd4,9'd4,9'd3,9'd2,-9'd4,9'd3,-9'd8,-9'd3,-9'd3,9'd8,9'd14,9'd24,9'd28,9'd35,9'd34,9'd31,9'd15,9'd8,-9'd5,-9'd5,-9'd18,-9'd24,-9'd16,-9'd13,-9'd1,-9'd4,-9'd4,-9'd3,9'd2,-9'd1,-9'd4,9'd1,9'd0,9'd2,-9'd3,-9'd5,-9'd1,-9'd12,-9'd6,-9'd6,-9'd8,-9'd6,9'd2,-9'd3,-9'd4,-9'd12,-9'd17,-9'd25,-9'd18,-9'd18,-9'd16,-9'd10,-9'd6,-9'd5,9'd2,-9'd2,9'd3,9'd3,-9'd3,-9'd3,-9'd2,9'd3,9'd0,-9'd3,-9'd2,-9'd5,-9'd11,-9'd24,-9'd25,-9'd26,-9'd26,-9'd31,-9'd30,-9'd24,-9'd23,-9'd18,-9'd17,-9'd13,-9'd3,-9'd1,9'd0,-9'd5,9'd2,9'd3,9'd1,-9'd2,9'd0,-9'd2,9'd4,9'd4,-9'd1,-9'd4,9'd1,9'd0,-9'd2,-9'd11,-9'd6,-9'd8,-9'd10,-9'd11,-9'd8,-9'd7,-9'd11,-9'd3,-9'd1,9'd1,9'd1,-9'd2,9'd2,9'd3,9'd2,-9'd3,-9'd2,9'd4,9'd3,9'd3,-9'd2,-9'd1,-9'd3,-9'd3,9'd3,-9'd4,-9'd1,9'd1,-9'd3,9'd1,-9'd2,9'd0,-9'd6,-9'd1,-9'd6,9'd2,9'd3,-9'd2,9'd0,-9'd3,-9'd3,-9'd2,-9'd2,9'd1,-9'd1,9'd0}; 
            // 1
            // weight_bin={-9'd4,-9'd3,-9'd4,-9'd3,9'd4,9'd2,-9'd4,-9'd1,9'd0,9'd2,9'd4,9'd1,9'd3,-9'd2,9'd0,-9'd3,9'd1,9'd4,9'd3,9'd5,-9'd2,-9'd1,9'd1,9'd4,-9'd4,-9'd2,9'd1,-9'd3,9'd2,9'd0,-9'd1,9'd2,9'd3,9'd4,9'd2,9'd0,9'd4,9'd4,-9'd2,9'd2,9'd1,-9'd2,-9'd1,-9'd1,-9'd3,-9'd2,9'd2,9'd3,9'd0,-9'd5,9'd2,-9'd1,9'd4,-9'd4,-9'd1,9'd4,9'd2,-9'd2,-9'd4,9'd0,9'd2,-9'd4,-9'd4,9'd0,-9'd1,9'd3,-9'd5,-9'd1,-9'd4,-9'd1,-9'd1,9'd4,-9'd5,-9'd6,-9'd5,-9'd7,9'd1,-9'd2,-9'd3,9'd3,-9'd1,9'd2,-9'd1,-9'd4,9'd1,9'd3,-9'd4,9'd0,9'd1,9'd0,9'd0,-9'd2,-9'd5,-9'd5,-9'd13,-9'd15,-9'd13,-9'd11,-9'd4,-9'd2,-9'd5,-9'd15,-9'd13,-9'd12,-9'd10,-9'd3,9'd1,9'd3,9'd2,9'd2,-9'd2,-9'd3,-9'd2,9'd4,-9'd1,9'd0,-9'd4,-9'd1,-9'd3,-9'd8,-9'd8,-9'd19,-9'd14,-9'd5,9'd4,9'd13,9'd9,9'd6,-9'd6,-9'd6,-9'd9,9'd4,9'd20,9'd24,9'd18,9'd6,9'd0,9'd1,-9'd4,9'd3,9'd1,-9'd4,9'd2,9'd3,9'd2,9'd1,-9'd5,-9'd14,-9'd24,-9'd28,-9'd25,-9'd1,9'd13,9'd13,9'd5,-9'd4,-9'd20,-9'd25,-9'd15,9'd2,9'd23,9'd33,9'd25,9'd10,-9'd3,-9'd3,9'd4,-9'd3,9'd0,9'd4,-9'd4,-9'd1,9'd4,-9'd3,-9'd10,-9'd23,-9'd37,-9'd53,-9'd45,-9'd21,-9'd2,-9'd2,-9'd15,-9'd41,-9'd42,-9'd46,-9'd25,-9'd6,9'd11,9'd16,9'd8,-9'd9,-9'd10,-9'd10,9'd2,9'd3,-9'd1,9'd2,9'd1,9'd3,-9'd4,-9'd8,-9'd20,-9'd24,-9'd51,-9'd62,-9'd57,-9'd36,-9'd19,-9'd25,-9'd36,-9'd38,-9'd48,-9'd45,-9'd29,9'd0,9'd1,-9'd5,-9'd12,-9'd25,-9'd21,-9'd8,9'd2,-9'd2,-9'd1,-9'd4,9'd3,9'd4,9'd3,-9'd8,-9'd20,-9'd33,-9'd48,-9'd66,-9'd69,-9'd53,-9'd34,-9'd15,-9'd12,-9'd5,-9'd20,-9'd17,-9'd12,-9'd14,-9'd25,-9'd27,-9'd42,-9'd40,-9'd24,-9'd11,9'd2,-9'd1,-9'd4,9'd1,-9'd3,9'd0,-9'd5,-9'd6,-9'd21,-9'd23,-9'd39,-9'd51,-9'd58,-9'd46,-9'd33,-9'd1,9'd27,9'd35,9'd19,-9'd9,-9'd16,-9'd31,-9'd38,-9'd49,-9'd52,-9'd35,-9'd21,-9'd6,-9'd5,9'd0,-9'd4,9'd0,9'd0,-9'd4,-9'd6,-9'd8,-9'd10,-9'd16,-9'd31,-9'd38,-9'd47,-9'd50,-9'd35,9'd15,9'd72,9'd81,9'd38,-9'd11,-9'd25,-9'd35,-9'd41,-9'd41,-9'd35,-9'd24,-9'd11,9'd2,9'd2,9'd1,-9'd3,-9'd3,9'd4,-9'd1,-9'd6,-9'd4,-9'd10,-9'd14,-9'd20,-9'd30,-9'd51,-9'd62,-9'd46,9'd27,9'd101,9'd101,9'd34,-9'd17,-9'd30,-9'd34,-9'd39,-9'd24,-9'd16,-9'd5,-9'd7,-9'd5,-9'd1,9'd1,9'd3,9'd4,9'd3,9'd1,-9'd2,-9'd3,-9'd9,-9'd10,-9'd23,-9'd33,-9'd62,-9'd79,-9'd46,9'd40,9'd110,9'd83,9'd10,-9'd22,-9'd33,-9'd36,-9'd33,-9'd13,-9'd7,-9'd6,-9'd2,-9'd1,-9'd3,-9'd2,9'd0,-9'd4,-9'd4,9'd1,-9'd3,-9'd4,-9'd5,-9'd14,-9'd18,-9'd46,-9'd81,-9'd89,-9'd42,9'd49,9'd110,9'd63,-9'd6,-9'd24,-9'd47,-9'd36,-9'd28,-9'd19,-9'd9,-9'd9,-9'd1,-9'd2,9'd0,-9'd2,9'd2,9'd4,-9'd1,-9'd3,-9'd5,9'd2,-9'd4,-9'd11,-9'd26,-9'd52,-9'd79,-9'd74,-9'd16,9'd60,9'd95,9'd54,-9'd13,-9'd56,-9'd51,-9'd36,-9'd22,-9'd18,-9'd11,-9'd4,-9'd2,9'd4,9'd2,9'd1,9'd1,-9'd4,-9'd2,9'd1,-9'd4,-9'd7,-9'd6,-9'd15,-9'd33,-9'd53,-9'd66,-9'd39,9'd10,9'd62,9'd85,9'd23,-9'd31,-9'd73,-9'd59,-9'd40,-9'd27,-9'd21,-9'd14,-9'd9,-9'd7,-9'd4,9'd3,9'd3,9'd4,-9'd3,9'd3,-9'd2,-9'd2,-9'd6,-9'd14,-9'd25,-9'd36,-9'd48,-9'd35,-9'd24,9'd8,9'd66,9'd75,9'd4,-9'd57,-9'd77,-9'd58,-9'd40,-9'd24,-9'd20,-9'd11,-9'd8,-9'd8,-9'd2,9'd3,9'd1,9'd1,9'd0,-9'd2,-9'd3,9'd3,-9'd10,-9'd21,-9'd32,-9'd37,-9'd30,-9'd13,-9'd7,9'd31,9'd71,9'd53,-9'd22,-9'd65,-9'd77,-9'd56,-9'd38,-9'd23,-9'd17,-9'd13,-9'd12,-9'd7,-9'd3,9'd3,9'd1,9'd0,9'd1,9'd3,9'd0,-9'd1,-9'd19,-9'd38,-9'd38,-9'd30,-9'd11,9'd2,9'd9,9'd33,9'd53,9'd37,-9'd29,-9'd54,-9'd50,-9'd49,-9'd31,-9'd24,-9'd17,-9'd21,-9'd19,-9'd10,9'd0,9'd0,9'd0,9'd0,9'd2,9'd0,-9'd5,-9'd10,-9'd23,-9'd43,-9'd31,-9'd18,-9'd1,-9'd6,9'd1,9'd17,9'd25,9'd7,-9'd23,-9'd35,-9'd31,-9'd39,-9'd27,-9'd27,-9'd25,-9'd24,-9'd12,-9'd10,9'd2,-9'd4,-9'd1,-9'd3,-9'd3,-9'd3,-9'd2,-9'd6,-9'd17,-9'd23,-9'd23,-9'd13,-9'd6,-9'd5,-9'd6,-9'd10,-9'd2,-9'd9,-9'd18,-9'd11,-9'd14,-9'd30,-9'd31,-9'd27,-9'd28,-9'd17,-9'd9,-9'd1,-9'd2,-9'd3,-9'd2,-9'd3,9'd0,9'd4,9'd4,9'd0,-9'd3,9'd1,9'd3,9'd5,-9'd9,-9'd17,-9'd23,-9'd36,-9'd35,-9'd22,-9'd1,9'd12,9'd2,-9'd15,-9'd31,-9'd29,-9'd19,-9'd20,-9'd6,-9'd8,-9'd3,-9'd1,9'd0,-9'd1,-9'd2,-9'd2,-9'd3,-9'd2,9'd13,9'd24,9'd18,9'd8,-9'd2,-9'd27,-9'd45,-9'd66,-9'd55,-9'd18,9'd10,9'd34,9'd34,9'd8,-9'd20,-9'd18,-9'd19,-9'd10,-9'd4,-9'd1,9'd1,9'd0,9'd3,9'd1,9'd4,9'd1,-9'd3,9'd7,9'd16,9'd31,9'd21,9'd14,-9'd9,-9'd20,-9'd39,-9'd40,-9'd34,-9'd14,9'd11,9'd38,9'd43,9'd6,-9'd6,-9'd13,-9'd12,-9'd6,9'd0,9'd2,9'd0,-9'd1,9'd0,9'd2,-9'd4,-9'd1,-9'd5,9'd1,9'd4,9'd9,9'd2,-9'd25,-9'd35,-9'd44,-9'd50,-9'd45,-9'd42,-9'd33,-9'd20,-9'd5,9'd0,9'd2,-9'd5,-9'd2,-9'd4,-9'd5,9'd0,-9'd2,9'd3,9'd4,-9'd5,9'd0,-9'd1,-9'd3,-9'd3,-9'd2,9'd1,-9'd1,-9'd7,-9'd15,-9'd18,-9'd28,-9'd30,-9'd29,-9'd35,-9'd25,-9'd26,-9'd18,-9'd7,-9'd3,-9'd4,9'd0,9'd0,-9'd1,9'd4,9'd3,9'd1,-9'd2,9'd1,-9'd3,9'd3,9'd4,-9'd1,9'd3,9'd4,-9'd1,-9'd3,-9'd2,-9'd2,-9'd8,-9'd5,-9'd7,-9'd4,-9'd7,-9'd1,9'd2,-9'd2,9'd1,-9'd1,-9'd2,-9'd3,9'd0,9'd1,-9'd1,9'd1,9'd3,9'd2,9'd2,9'd1,-9'd4,-9'd3,-9'd3,9'd3,-9'd4,-9'd4,9'd3,9'd3,-9'd4,9'd3,-9'd1,9'd1,-9'd3,-9'd1,9'd1,9'd3,9'd3,-9'd2,-9'd3,9'd0,9'd1,9'd3,-9'd5,9'd0,9'd0,-9'd2};
            // 2
            // weight_bin={9'd4,-9'd1,-9'd4,-9'd3,9'd0,-9'd3,9'd1,9'd4,9'd0,-9'd1,9'd4,9'd3,9'd3,9'd0,9'd0,-9'd4,9'd0,9'd4,9'd0,-9'd4,9'd3,9'd4,9'd4,9'd0,9'd1,9'd1,-9'd2,-9'd1,9'd4,9'd0,9'd4,-9'd3,-9'd1,9'd0,-9'd3,9'd3,9'd3,-9'd3,9'd4,9'd4,-9'd3,9'd0,9'd5,-9'd3,9'd1,-9'd3,9'd3,9'd0,9'd1,9'd3,-9'd1,-9'd5,9'd0,9'd0,9'd2,9'd2,-9'd2,-9'd2,9'd3,9'd1,9'd1,9'd2,9'd2,-9'd3,9'd0,9'd0,-9'd5,9'd4,9'd5,9'd8,-9'd1,9'd9,9'd4,9'd5,-9'd1,-9'd5,-9'd6,-9'd5,-9'd6,9'd0,9'd2,9'd1,-9'd3,9'd2,9'd4,-9'd1,9'd2,9'd0,9'd2,-9'd3,-9'd3,9'd3,9'd3,9'd20,9'd27,9'd29,9'd32,9'd33,9'd19,9'd12,9'd14,9'd7,-9'd7,-9'd8,-9'd13,-9'd11,-9'd9,-9'd7,9'd2,9'd3,-9'd2,-9'd1,-9'd1,9'd0,9'd1,9'd4,-9'd5,9'd3,9'd1,9'd8,9'd28,9'd39,9'd47,9'd54,9'd51,9'd41,9'd36,9'd25,9'd29,9'd19,9'd6,-9'd2,-9'd22,-9'd23,-9'd20,-9'd16,-9'd8,9'd1,9'd4,-9'd1,9'd0,9'd2,9'd1,9'd1,9'd2,9'd5,9'd9,9'd23,9'd40,9'd50,9'd55,9'd56,9'd50,9'd55,9'd56,9'd50,9'd49,9'd35,9'd17,-9'd9,-9'd18,-9'd26,-9'd28,-9'd18,-9'd10,-9'd2,9'd2,-9'd1,9'd1,-9'd5,9'd3,-9'd5,-9'd1,-9'd2,9'd14,9'd35,9'd32,9'd35,9'd36,9'd25,9'd19,9'd25,9'd25,9'd22,9'd20,9'd6,9'd3,-9'd12,-9'd18,-9'd20,-9'd29,-9'd26,-9'd9,-9'd5,-9'd3,9'd4,-9'd2,-9'd4,-9'd3,9'd0,9'd0,9'd10,9'd26,9'd30,9'd24,9'd19,9'd9,9'd8,9'd8,9'd10,9'd16,9'd7,-9'd3,-9'd21,-9'd10,-9'd3,-9'd12,-9'd16,-9'd17,-9'd29,-9'd16,-9'd5,-9'd2,9'd4,-9'd2,9'd4,9'd0,9'd1,9'd1,9'd13,9'd19,9'd11,9'd13,9'd8,9'd6,9'd15,9'd7,9'd15,9'd28,9'd20,-9'd3,-9'd8,-9'd5,9'd0,-9'd11,-9'd14,-9'd12,-9'd33,-9'd25,-9'd5,9'd4,9'd1,-9'd3,9'd1,-9'd3,9'd2,9'd4,9'd12,-9'd3,-9'd13,-9'd23,-9'd23,-9'd7,-9'd12,-9'd20,-9'd13,9'd1,9'd10,9'd7,-9'd2,-9'd6,-9'd8,-9'd15,-9'd15,-9'd18,-9'd32,-9'd21,-9'd1,-9'd4,-9'd2,-9'd4,9'd3,9'd4,-9'd4,-9'd1,-9'd8,-9'd30,-9'd53,-9'd59,-9'd52,-9'd46,-9'd65,-9'd73,-9'd79,-9'd50,-9'd19,-9'd2,-9'd7,-9'd9,-9'd13,-9'd11,-9'd15,-9'd21,-9'd28,-9'd13,-9'd2,-9'd2,9'd3,9'd4,9'd1,9'd4,-9'd4,-9'd6,-9'd30,-9'd70,-9'd98,-9'd102,-9'd100,-9'd106,-9'd109,-9'd120,-9'd127,-9'd93,-9'd47,-9'd24,-9'd17,-9'd16,-9'd1,-9'd12,-9'd14,-9'd29,-9'd22,-9'd7,9'd1,9'd2,9'd4,-9'd3,9'd1,-9'd4,-9'd1,-9'd16,-9'd50,-9'd102,-9'd120,-9'd119,-9'd117,-9'd122,-9'd115,-9'd120,-9'd118,-9'd96,-9'd57,-9'd46,-9'd45,-9'd22,-9'd4,-9'd6,-9'd17,-9'd36,-9'd31,-9'd13,-9'd1,-9'd5,-9'd1,-9'd1,9'd2,-9'd1,9'd1,-9'd12,-9'd59,-9'd101,-9'd110,-9'd102,-9'd83,-9'd75,-9'd62,-9'd60,-9'd54,-9'd56,-9'd51,-9'd41,-9'd43,-9'd31,-9'd13,-9'd17,-9'd22,-9'd38,-9'd32,-9'd15,9'd7,9'd4,9'd5,9'd1,9'd3,-9'd4,-9'd4,-9'd8,-9'd45,-9'd63,-9'd51,-9'd34,-9'd21,-9'd13,-9'd1,9'd8,9'd11,-9'd11,-9'd23,-9'd22,-9'd32,-9'd23,-9'd24,-9'd27,-9'd33,-9'd35,-9'd35,-9'd14,9'd1,9'd9,9'd4,9'd5,9'd4,-9'd1,9'd3,9'd5,-9'd11,-9'd16,-9'd2,9'd4,9'd15,9'd17,9'd17,9'd22,9'd23,9'd5,-9'd7,-9'd10,-9'd25,-9'd36,-9'd23,-9'd29,-9'd25,-9'd24,-9'd21,9'd1,9'd9,9'd8,-9'd2,9'd0,-9'd3,9'd0,-9'd1,9'd16,9'd22,9'd26,9'd22,9'd16,9'd17,9'd13,9'd21,9'd30,9'd21,9'd1,9'd1,-9'd5,-9'd19,-9'd21,-9'd19,-9'd13,-9'd3,9'd3,9'd2,9'd14,9'd25,9'd8,-9'd1,9'd2,-9'd4,-9'd7,9'd1,9'd26,9'd51,9'd49,9'd31,9'd23,9'd19,9'd30,9'd31,9'd41,9'd26,9'd13,9'd18,9'd7,9'd0,-9'd7,-9'd1,9'd7,9'd11,9'd19,9'd29,9'd40,9'd34,9'd14,9'd2,-9'd4,9'd4,-9'd7,9'd7,9'd36,9'd58,9'd50,9'd42,9'd23,9'd32,9'd44,9'd53,9'd59,9'd54,9'd34,9'd15,9'd13,9'd10,9'd6,9'd6,9'd16,9'd23,9'd32,9'd51,9'd66,9'd34,9'd2,-9'd1,-9'd1,9'd2,-9'd1,9'd5,9'd20,9'd37,9'd50,9'd45,9'd45,9'd45,9'd45,9'd47,9'd49,9'd29,9'd18,9'd2,9'd8,9'd13,9'd15,9'd13,9'd19,9'd32,9'd52,9'd61,9'd52,9'd26,9'd7,-9'd1,-9'd2,-9'd4,-9'd6,9'd1,9'd19,9'd29,9'd40,9'd44,9'd42,9'd32,9'd35,9'd31,9'd13,9'd0,9'd3,-9'd4,9'd2,9'd11,9'd20,9'd35,9'd30,9'd44,9'd59,9'd60,9'd39,9'd14,9'd6,9'd3,9'd4,9'd4,9'd4,9'd0,9'd10,9'd14,9'd18,9'd26,9'd32,9'd32,9'd22,9'd15,-9'd10,-9'd18,-9'd13,9'd0,9'd8,9'd15,9'd28,9'd31,9'd31,9'd48,9'd51,9'd55,9'd25,9'd5,9'd2,9'd3,9'd0,-9'd4,9'd0,9'd0,9'd8,9'd7,9'd8,9'd13,9'd14,9'd12,9'd10,9'd1,-9'd12,-9'd28,-9'd31,-9'd25,-9'd17,9'd0,9'd22,9'd25,9'd37,9'd35,9'd31,9'd24,9'd16,9'd7,9'd1,9'd0,9'd4,9'd3,9'd3,-9'd3,9'd1,-9'd2,-9'd19,-9'd17,-9'd31,-9'd24,-9'd16,-9'd16,-9'd27,-9'd48,-9'd50,-9'd52,-9'd38,-9'd33,-9'd4,9'd5,9'd8,9'd22,9'd13,9'd8,9'd4,-9'd2,-9'd4,-9'd2,9'd1,9'd4,9'd0,-9'd2,-9'd7,-9'd13,-9'd18,-9'd30,-9'd38,-9'd47,-9'd45,-9'd38,-9'd34,-9'd41,-9'd40,-9'd40,-9'd36,-9'd31,-9'd21,-9'd20,-9'd13,-9'd8,-9'd6,-9'd4,9'd1,9'd5,9'd1,9'd0,-9'd3,-9'd2,-9'd1,-9'd4,-9'd1,-9'd2,-9'd7,-9'd19,-9'd24,-9'd19,-9'd23,-9'd24,-9'd19,-9'd18,-9'd21,-9'd19,-9'd20,-9'd10,-9'd11,-9'd6,-9'd2,-9'd7,-9'd5,-9'd2,9'd0,9'd3,9'd0,9'd1,-9'd1,9'd2,9'd1,-9'd4,9'd2,-9'd1,9'd3,-9'd6,-9'd2,9'd0,9'd1,-9'd2,-9'd4,-9'd5,-9'd5,9'd2,-9'd5,-9'd3,9'd1,9'd2,-9'd5,9'd1,9'd0,9'd4,9'd0,9'd2,9'd0,9'd4,9'd0,-9'd3,9'd1,-9'd2,9'd1,9'd3,-9'd4,-9'd3,9'd0,9'd0,-9'd2,9'd4,9'd2,-9'd2,9'd0,-9'd1,-9'd3,9'd2,-9'd3,9'd1,9'd3,-9'd4,9'd0,9'd4,9'd2,-9'd2,9'd1,-9'd4};
            // 3 
            // weight_bin={9'd1,9'd4,9'd4,9'd0,9'd2,-9'd1,-9'd1,9'd0,-9'd3,9'd2,9'd2,-9'd1,-9'd1,-9'd3,9'd1,9'd2,9'd4,-9'd4,-9'd4,9'd0,9'd4,9'd0,9'd1,9'd1,-9'd1,9'd3,9'd3,-9'd3,-9'd3,-9'd4,-9'd1,9'd0,9'd4,-9'd4,9'd3,-9'd3,9'd0,9'd0,9'd3,-9'd4,-9'd3,9'd0,9'd2,-9'd2,9'd1,-9'd1,-9'd4,9'd0,-9'd1,9'd3,9'd3,9'd3,9'd3,-9'd4,-9'd4,9'd1,9'd1,-9'd4,9'd4,9'd0,-9'd3,9'd3,9'd4,9'd1,-9'd2,9'd0,-9'd4,9'd2,9'd2,-9'd2,-9'd5,9'd2,-9'd5,-9'd4,9'd2,-9'd3,9'd0,9'd3,-9'd1,-9'd1,9'd4,9'd1,9'd2,-9'd2,-9'd4,9'd1,-9'd3,-9'd2,-9'd4,9'd4,-9'd3,9'd2,9'd2,9'd7,9'd10,9'd10,9'd25,9'd21,9'd23,9'd17,9'd9,9'd12,9'd2,9'd1,-9'd1,-9'd7,-9'd5,-9'd5,-9'd2,-9'd3,9'd0,9'd1,9'd4,9'd1,-9'd1,-9'd2,9'd2,9'd10,9'd6,9'd11,9'd26,9'd24,9'd33,9'd34,9'd35,9'd35,9'd27,9'd16,9'd4,-9'd1,-9'd4,-9'd7,-9'd24,-9'd23,-9'd18,-9'd18,-9'd4,9'd3,-9'd2,9'd4,9'd0,-9'd1,9'd2,9'd4,9'd12,9'd23,9'd24,9'd28,9'd33,9'd29,9'd33,9'd27,9'd22,9'd20,9'd7,9'd14,9'd9,-9'd8,-9'd13,-9'd18,-9'd30,-9'd34,-9'd40,-9'd35,-9'd10,-9'd4,9'd3,9'd2,-9'd2,-9'd1,-9'd2,9'd6,9'd18,9'd31,9'd32,9'd27,9'd32,9'd31,9'd27,9'd22,9'd26,9'd34,9'd29,9'd20,9'd25,9'd17,9'd11,-9'd7,-9'd4,-9'd24,-9'd41,-9'd41,-9'd16,-9'd6,-9'd1,9'd4,9'd2,-9'd4,9'd3,9'd7,9'd29,9'd39,9'd37,9'd25,9'd10,9'd8,9'd11,9'd6,9'd15,9'd17,9'd31,9'd25,9'd13,9'd14,9'd8,9'd11,9'd14,-9'd4,-9'd25,-9'd39,-9'd32,-9'd4,9'd2,-9'd4,-9'd1,9'd3,-9'd3,9'd14,9'd32,9'd34,9'd28,9'd4,9'd1,-9'd8,9'd0,-9'd16,-9'd13,9'd0,9'd29,9'd40,9'd25,9'd17,9'd17,9'd21,9'd23,9'd7,-9'd19,-9'd47,-9'd29,-9'd9,9'd1,9'd1,9'd2,9'd0,-9'd1,9'd12,9'd22,9'd13,9'd7,-9'd10,-9'd31,-9'd42,-9'd64,-9'd87,-9'd70,-9'd29,9'd30,9'd58,9'd40,9'd23,9'd23,9'd19,9'd33,9'd14,-9'd19,-9'd41,-9'd21,-9'd6,9'd4,9'd4,9'd0,9'd1,-9'd2,9'd5,9'd6,9'd2,-9'd22,-9'd54,-9'd80,-9'd101,-9'd116,-9'd116,-9'd85,-9'd26,9'd37,9'd49,9'd39,9'd31,9'd28,9'd26,9'd31,9'd2,-9'd15,-9'd20,-9'd13,-9'd5,9'd4,9'd4,9'd4,9'd2,9'd2,9'd8,9'd2,-9'd23,-9'd53,-9'd81,-9'd100,-9'd88,-9'd78,-9'd53,-9'd33,9'd1,9'd29,9'd31,9'd29,9'd28,9'd25,9'd22,9'd9,-9'd10,-9'd15,-9'd17,-9'd2,-9'd2,9'd1,-9'd2,9'd4,-9'd1,9'd0,-9'd4,-9'd4,-9'd33,-9'd54,-9'd71,-9'd63,-9'd44,-9'd32,-9'd18,-9'd2,9'd14,9'd41,9'd25,9'd25,9'd17,9'd6,-9'd16,-9'd26,-9'd31,-9'd25,-9'd18,-9'd3,-9'd4,9'd1,-9'd4,9'd1,9'd2,-9'd4,-9'd1,-9'd11,-9'd23,-9'd46,-9'd52,-9'd43,-9'd27,-9'd24,-9'd15,9'd10,9'd29,9'd29,9'd7,9'd9,9'd7,-9'd8,-9'd29,-9'd41,-9'd33,-9'd34,-9'd17,-9'd4,9'd1,9'd2,9'd1,-9'd4,-9'd1,9'd3,9'd0,-9'd2,-9'd17,-9'd39,-9'd47,-9'd35,-9'd27,-9'd39,-9'd22,9'd10,9'd16,9'd5,-9'd12,-9'd14,-9'd10,9'd1,-9'd12,-9'd13,-9'd20,-9'd22,-9'd9,-9'd3,9'd3,9'd1,-9'd4,-9'd3,9'd3,-9'd4,9'd6,-9'd2,-9'd16,-9'd31,-9'd46,-9'd48,-9'd43,-9'd39,-9'd19,9'd4,9'd15,-9'd5,-9'd24,-9'd27,-9'd11,9'd5,9'd11,9'd12,9'd11,-9'd7,-9'd9,-9'd3,9'd2,-9'd2,-9'd4,9'd1,9'd0,9'd4,9'd5,9'd7,-9'd5,-9'd21,-9'd37,-9'd65,-9'd80,-9'd77,-9'd49,-9'd24,-9'd11,-9'd29,-9'd43,-9'd23,-9'd8,9'd15,9'd24,9'd23,9'd25,9'd15,-9'd1,-9'd1,-9'd5,9'd3,9'd0,9'd0,9'd0,9'd3,9'd17,9'd9,9'd1,-9'd22,-9'd42,-9'd71,-9'd115,-9'd127,-9'd119,-9'd100,-9'd80,-9'd77,-9'd44,-9'd10,9'd6,9'd18,9'd37,9'd16,9'd32,9'd23,9'd2,-9'd14,-9'd8,-9'd3,9'd0,9'd2,9'd2,9'd8,9'd32,9'd29,9'd20,-9'd8,-9'd22,-9'd52,-9'd93,-9'd117,-9'd120,-9'd122,-9'd120,-9'd87,-9'd34,9'd13,9'd16,9'd31,9'd39,9'd30,9'd35,9'd24,9'd0,-9'd10,-9'd8,-9'd2,9'd0,9'd4,9'd4,9'd4,9'd32,9'd45,9'd33,9'd16,9'd6,-9'd14,-9'd37,-9'd48,-9'd63,-9'd76,-9'd74,-9'd46,-9'd15,9'd22,9'd27,9'd40,9'd39,9'd36,9'd32,9'd7,-9'd6,-9'd7,-9'd7,9'd3,-9'd2,9'd1,-9'd2,9'd8,9'd31,9'd44,9'd41,9'd36,9'd21,9'd12,9'd7,-9'd3,-9'd21,-9'd27,-9'd21,-9'd12,9'd0,9'd19,9'd29,9'd31,9'd23,9'd30,9'd13,-9'd8,-9'd14,-9'd8,9'd2,9'd1,9'd1,-9'd2,-9'd1,9'd7,9'd27,9'd42,9'd41,9'd33,9'd25,9'd21,9'd16,9'd8,-9'd7,-9'd1,-9'd4,-9'd2,-9'd2,9'd10,9'd14,9'd24,9'd27,9'd16,-9'd10,-9'd18,-9'd18,-9'd3,-9'd2,-9'd5,-9'd2,-9'd3,9'd1,9'd3,9'd16,9'd33,9'd34,9'd36,9'd26,9'd15,9'd17,9'd17,9'd14,-9'd1,-9'd7,-9'd1,-9'd2,9'd6,9'd5,9'd4,9'd10,9'd0,-9'd17,-9'd13,-9'd11,-9'd1,9'd3,-9'd4,-9'd3,9'd4,9'd4,9'd3,9'd7,9'd25,9'd32,9'd38,9'd36,9'd17,9'd23,9'd8,9'd8,9'd2,9'd7,9'd1,9'd3,-9'd4,-9'd1,9'd7,-9'd4,-9'd10,-9'd16,-9'd12,-9'd4,-9'd1,-9'd1,9'd2,9'd2,-9'd1,9'd0,9'd0,9'd4,9'd10,9'd21,9'd27,9'd40,9'd34,9'd27,9'd41,9'd37,9'd30,9'd27,9'd25,9'd9,-9'd1,-9'd7,-9'd17,-9'd16,-9'd16,-9'd10,-9'd6,9'd1,9'd3,9'd0,-9'd2,9'd4,9'd0,-9'd3,9'd3,9'd5,9'd6,9'd9,9'd13,9'd5,9'd16,9'd19,9'd21,9'd31,9'd27,9'd21,9'd15,9'd0,-9'd10,-9'd18,-9'd14,-9'd14,-9'd6,-9'd10,-9'd4,9'd1,9'd0,9'd3,9'd2,9'd0,9'd1,9'd3,-9'd4,-9'd2,9'd3,-9'd4,9'd2,9'd2,9'd0,-9'd5,-9'd5,-9'd3,-9'd5,-9'd3,-9'd4,-9'd4,-9'd1,-9'd9,-9'd8,9'd0,-9'd4,-9'd5,-9'd2,9'd3,-9'd1,9'd2,9'd3,-9'd1,9'd2,9'd1,-9'd3,-9'd1,9'd3,9'd2,9'd1,-9'd1,-9'd3,-9'd2,9'd3,9'd0,-9'd3,9'd0,-9'd4,-9'd1,-9'd1,-9'd5,-9'd3,-9'd3,-9'd3,9'd4,9'd2,-9'd3,-9'd2,9'd3,9'd4,9'd0};
            // 4 
            // weight_bin={9'd0,-9'd3,9'd3,-9'd1,9'd0,-9'd1,9'd2,9'd1,-9'd1,-9'd1,9'd0,-9'd4,9'd0,-9'd4,9'd4,9'd2,9'd0,9'd3,9'd0,9'd4,9'd1,9'd2,9'd1,-9'd3,-9'd4,-9'd2,9'd4,9'd2,-9'd1,-9'd3,9'd5,9'd0,-9'd4,-9'd2,9'd0,-9'd2,-9'd3,9'd0,-9'd6,-9'd1,-9'd9,9'd0,9'd3,9'd3,-9'd7,-9'd2,-9'd1,-9'd4,9'd2,-9'd2,9'd0,9'd2,-9'd4,9'd1,-9'd2,9'd3,9'd4,-9'd1,-9'd3,9'd3,-9'd3,9'd4,9'd3,-9'd1,-9'd7,-9'd3,-9'd8,-9'd14,-9'd22,-9'd19,-9'd15,-9'd12,-9'd17,-9'd4,-9'd7,-9'd1,-9'd3,-9'd4,-9'd2,9'd0,-9'd4,-9'd2,9'd3,9'd0,-9'd2,9'd4,-9'd4,-9'd1,9'd4,9'd0,-9'd3,-9'd9,-9'd13,-9'd19,-9'd23,-9'd26,-9'd35,-9'd47,-9'd41,-9'd40,-9'd31,-9'd19,-9'd11,-9'd9,-9'd2,9'd1,-9'd2,9'd2,-9'd4,9'd3,-9'd4,9'd2,-9'd4,-9'd1,9'd0,-9'd1,9'd0,-9'd3,-9'd6,-9'd5,-9'd12,-9'd21,-9'd35,-9'd37,-9'd46,-9'd53,-9'd54,-9'd43,-9'd27,-9'd30,-9'd20,-9'd5,9'd3,-9'd2,9'd3,9'd3,9'd3,-9'd4,9'd1,9'd3,9'd3,-9'd4,-9'd1,9'd2,9'd3,9'd5,9'd5,-9'd1,-9'd3,-9'd4,-9'd22,-9'd30,-9'd40,-9'd44,-9'd34,-9'd17,-9'd7,-9'd4,-9'd4,9'd8,9'd12,9'd15,9'd26,9'd34,9'd14,9'd5,-9'd3,9'd4,9'd0,-9'd3,9'd0,-9'd2,9'd4,9'd9,9'd3,9'd7,9'd0,-9'd10,-9'd21,-9'd44,-9'd66,-9'd69,-9'd86,-9'd73,-9'd55,-9'd45,-9'd42,-9'd19,-9'd8,9'd15,9'd43,9'd50,9'd17,9'd4,-9'd4,-9'd2,9'd4,9'd2,9'd0,-9'd2,-9'd1,9'd8,9'd2,9'd1,-9'd13,-9'd23,-9'd37,-9'd60,-9'd76,-9'd71,-9'd95,-9'd109,-9'd88,-9'd64,-9'd53,-9'd33,-9'd25,-9'd1,9'd28,9'd33,9'd8,9'd3,-9'd2,-9'd4,-9'd3,-9'd3,-9'd5,9'd2,9'd4,-9'd1,-9'd1,-9'd3,-9'd22,-9'd18,-9'd34,-9'd44,-9'd52,-9'd54,-9'd97,-9'd109,-9'd81,-9'd47,-9'd38,-9'd21,-9'd15,-9'd10,9'd11,9'd7,-9'd10,-9'd15,-9'd1,-9'd1,9'd2,-9'd3,-9'd1,-9'd1,-9'd2,9'd2,-9'd12,-9'd12,-9'd17,-9'd17,-9'd18,-9'd19,-9'd21,-9'd43,-9'd116,-9'd99,-9'd38,-9'd25,-9'd20,-9'd13,-9'd21,-9'd19,-9'd8,-9'd10,-9'd17,-9'd14,-9'd7,9'd2,-9'd1,9'd1,9'd1,-9'd4,9'd1,-9'd4,-9'd22,-9'd14,-9'd6,9'd9,9'd7,9'd3,9'd6,-9'd41,-9'd107,-9'd58,9'd3,9'd5,-9'd9,-9'd4,-9'd22,-9'd17,-9'd11,-9'd17,-9'd11,-9'd5,-9'd3,9'd1,9'd3,9'd2,-9'd3,9'd0,-9'd6,-9'd10,-9'd9,-9'd5,9'd11,9'd29,9'd37,9'd38,9'd28,-9'd51,-9'd87,-9'd14,9'd33,9'd21,-9'd2,-9'd9,-9'd30,-9'd20,-9'd17,-9'd21,-9'd11,-9'd5,-9'd3,-9'd1,9'd0,-9'd2,-9'd5,9'd2,-9'd3,-9'd6,9'd7,9'd25,9'd37,9'd39,9'd60,9'd85,9'd58,-9'd18,-9'd53,9'd11,9'd45,9'd19,-9'd1,-9'd14,-9'd18,-9'd10,-9'd12,-9'd16,-9'd12,-9'd1,9'd2,9'd4,9'd4,-9'd4,-9'd3,9'd0,9'd3,9'd19,9'd41,9'd48,9'd61,9'd53,9'd79,9'd104,9'd70,-9'd9,-9'd19,9'd19,9'd45,9'd36,9'd19,9'd9,9'd10,9'd6,9'd3,-9'd9,-9'd7,-9'd2,9'd3,-9'd4,-9'd4,9'd4,-9'd1,-9'd4,9'd17,9'd29,9'd56,9'd66,9'd55,9'd45,9'd66,9'd69,9'd47,9'd9,-9'd9,9'd14,9'd47,9'd60,9'd41,9'd39,9'd20,9'd16,9'd11,9'd1,9'd2,-9'd2,9'd4,9'd3,9'd1,9'd2,9'd0,9'd1,9'd11,9'd23,9'd40,9'd51,9'd51,9'd42,9'd32,9'd27,9'd21,9'd5,9'd6,9'd38,9'd69,9'd65,9'd44,9'd29,9'd2,9'd4,9'd4,9'd2,-9'd7,9'd2,-9'd2,-9'd1,-9'd4,-9'd2,9'd0,9'd1,9'd5,9'd12,9'd27,9'd45,9'd54,9'd34,9'd8,9'd2,9'd13,9'd20,9'd46,9'd69,9'd72,9'd55,9'd27,9'd9,9'd11,9'd9,-9'd2,-9'd3,-9'd7,9'd0,9'd0,-9'd2,9'd4,9'd4,-9'd3,-9'd4,-9'd8,-9'd14,9'd8,9'd28,9'd49,9'd34,9'd8,9'd6,9'd12,9'd42,9'd63,9'd65,9'd53,9'd22,9'd2,-9'd19,-9'd7,-9'd12,-9'd21,-9'd19,-9'd13,-9'd3,9'd0,9'd0,-9'd2,-9'd4,9'd3,-9'd9,-9'd13,-9'd26,-9'd19,-9'd9,-9'd2,-9'd2,-9'd22,-9'd27,-9'd8,9'd15,9'd33,9'd32,9'd10,-9'd19,-9'd32,-9'd39,-9'd34,-9'd28,-9'd39,-9'd22,-9'd15,-9'd4,-9'd5,9'd2,-9'd3,-9'd4,-9'd2,-9'd2,-9'd16,-9'd35,-9'd46,-9'd59,-9'd66,-9'd74,-9'd75,-9'd68,-9'd62,-9'd26,-9'd7,-9'd8,-9'd18,-9'd27,-9'd31,-9'd37,-9'd36,-9'd37,-9'd36,-9'd21,-9'd11,9'd1,9'd4,9'd4,9'd4,-9'd4,-9'd2,-9'd2,-9'd14,-9'd33,-9'd56,-9'd73,-9'd86,-9'd91,-9'd86,-9'd72,-9'd56,-9'd51,-9'd25,-9'd14,-9'd20,-9'd11,-9'd21,-9'd33,-9'd30,-9'd23,-9'd26,-9'd17,-9'd8,-9'd6,9'd0,9'd1,-9'd1,-9'd3,-9'd3,9'd1,-9'd4,-9'd25,-9'd46,-9'd60,-9'd66,-9'd69,-9'd65,-9'd44,-9'd37,-9'd35,-9'd33,-9'd18,-9'd21,-9'd3,-9'd8,-9'd10,-9'd8,-9'd15,-9'd11,-9'd7,-9'd6,-9'd3,9'd1,9'd0,9'd1,9'd0,-9'd1,-9'd2,-9'd2,-9'd15,-9'd26,-9'd30,-9'd34,-9'd37,-9'd34,-9'd26,-9'd29,-9'd29,-9'd29,-9'd7,-9'd9,-9'd5,9'd14,9'd15,9'd14,9'd3,-9'd6,9'd1,-9'd3,-9'd2,-9'd2,9'd2,9'd2,-9'd2,-9'd3,9'd0,9'd1,-9'd3,-9'd15,-9'd15,-9'd22,-9'd21,-9'd20,-9'd18,-9'd21,-9'd24,-9'd17,-9'd13,-9'd1,9'd11,9'd23,9'd21,9'd14,9'd2,9'd1,9'd1,-9'd2,-9'd2,-9'd1,-9'd2,-9'd2,9'd4,-9'd2,9'd4,9'd3,-9'd4,-9'd3,-9'd15,-9'd11,-9'd18,-9'd17,-9'd13,-9'd19,-9'd27,-9'd30,-9'd22,-9'd20,-9'd10,-9'd5,9'd0,9'd1,-9'd7,-9'd6,-9'd5,9'd4,9'd2,-9'd4,-9'd1,9'd4,-9'd4,9'd0,-9'd3,-9'd4,-9'd3,-9'd5,-9'd19,-9'd22,-9'd33,-9'd35,-9'd47,-9'd47,-9'd46,-9'd43,-9'd50,-9'd48,-9'd60,-9'd48,-9'd29,-9'd27,-9'd14,-9'd5,-9'd1,9'd3,-9'd1,9'd3,-9'd3,-9'd4,-9'd3,9'd2,9'd0,-9'd1,-9'd1,-9'd5,-9'd5,-9'd11,-9'd20,-9'd26,-9'd35,-9'd32,-9'd35,-9'd47,-9'd35,-9'd33,-9'd28,-9'd26,-9'd18,-9'd6,-9'd2,9'd1,-9'd2,-9'd2,9'd0,9'd4,-9'd2,-9'd2,-9'd2,-9'd4,9'd2,-9'd1,9'd0,9'd4,9'd1,9'd3,9'd0,-9'd2,9'd2,-9'd1,-9'd4,-9'd5,-9'd4,-9'd2,9'd0,9'd1,9'd3,-9'd4,9'd0,9'd2,9'd3,-9'd3,-9'd4,9'd2,-9'd3};
            // 5
            //  weight_bin={9'd5,-9'd3,9'd2,-9'd1,-9'd4,-9'd4,9'd2,-9'd1,-9'd3,9'd5,9'd3,9'd3,-9'd2,9'd0,9'd1,-9'd1,9'd2,-9'd1,-9'd1,9'd0,-9'd2,-9'd3,-9'd1,-9'd2,-9'd1,-9'd2,9'd2,-9'd1,9'd4,9'd1,-9'd2,9'd5,-9'd1,-9'd4,9'd3,-9'd3,9'd3,9'd3,-9'd1,-9'd2,9'd2,9'd2,9'd4,9'd1,9'd0,9'd4,9'd1,-9'd4,-9'd1,9'd0,9'd2,-9'd4,-9'd5,-9'd3,9'd1,9'd3,-9'd4,9'd2,9'd0,9'd4,-9'd3,-9'd1,9'd1,-9'd4,9'd3,-9'd2,9'd1,-9'd3,9'd3,9'd0,-9'd1,-9'd4,-9'd5,-9'd1,-9'd5,-9'd1,9'd3,9'd0,-9'd2,-9'd2,9'd2,-9'd4,-9'd4,9'd0,9'd3,-9'd3,-9'd1,-9'd2,9'd3,-9'd2,-9'd1,9'd1,-9'd3,9'd0,-9'd10,-9'd12,-9'd9,-9'd12,-9'd12,-9'd10,-9'd12,-9'd2,-9'd6,-9'd8,-9'd4,-9'd4,-9'd7,-9'd3,-9'd7,-9'd3,9'd3,9'd2,9'd2,9'd2,-9'd2,-9'd4,9'd0,9'd0,-9'd2,-9'd10,-9'd20,-9'd25,-9'd28,-9'd33,-9'd33,-9'd38,-9'd24,-9'd13,9'd1,9'd6,-9'd5,-9'd5,-9'd10,9'd4,9'd7,9'd14,9'd7,-9'd1,9'd4,-9'd5,9'd4,9'd1,9'd3,9'd1,-9'd7,-9'd9,-9'd20,-9'd22,-9'd20,-9'd16,-9'd8,-9'd4,-9'd12,-9'd21,-9'd8,-9'd1,9'd6,9'd13,9'd17,9'd9,9'd16,9'd23,9'd29,9'd44,9'd32,9'd19,9'd7,9'd4,9'd1,-9'd2,-9'd3,-9'd7,-9'd10,-9'd21,-9'd22,-9'd26,-9'd11,9'd0,9'd13,9'd19,9'd5,9'd7,9'd2,-9'd4,-9'd8,9'd0,9'd10,9'd19,9'd18,9'd23,9'd51,9'd73,9'd66,9'd37,9'd17,9'd4,-9'd1,-9'd2,9'd1,-9'd3,-9'd25,-9'd28,-9'd26,-9'd15,9'd8,9'd11,9'd26,9'd20,9'd6,-9'd9,-9'd14,-9'd17,-9'd17,9'd0,9'd5,9'd18,9'd21,9'd32,9'd52,9'd79,9'd92,9'd61,9'd19,9'd1,-9'd4,-9'd3,-9'd3,-9'd12,-9'd31,-9'd33,-9'd26,-9'd8,9'd10,9'd13,9'd17,9'd17,9'd7,-9'd19,-9'd39,-9'd32,-9'd31,-9'd13,9'd1,9'd15,9'd34,9'd52,9'd65,9'd95,9'd121,9'd86,9'd19,9'd3,9'd3,9'd3,-9'd2,-9'd6,-9'd16,-9'd24,-9'd18,9'd3,9'd25,9'd21,9'd24,9'd43,9'd26,-9'd1,-9'd38,-9'd48,-9'd58,-9'd35,-9'd17,9'd2,9'd28,9'd42,9'd57,9'd86,9'd105,9'd81,9'd16,9'd6,9'd0,-9'd1,-9'd2,-9'd6,-9'd11,-9'd7,9'd0,9'd15,9'd36,9'd40,9'd45,9'd51,9'd55,9'd19,-9'd12,-9'd45,-9'd62,-9'd69,-9'd79,-9'd79,-9'd60,-9'd47,-9'd31,-9'd13,9'd18,9'd33,9'd2,-9'd2,9'd2,9'd2,-9'd2,-9'd7,9'd1,9'd6,9'd12,9'd32,9'd34,9'd31,9'd40,9'd54,9'd68,9'd40,-9'd15,-9'd53,-9'd69,-9'd78,-9'd94,-9'd124,-9'd127,-9'd127,-9'd105,-9'd76,-9'd31,-9'd1,9'd0,-9'd1,-9'd4,-9'd2,-9'd2,9'd4,-9'd1,9'd8,9'd16,9'd23,9'd25,9'd10,9'd41,9'd74,9'd79,9'd50,-9'd12,-9'd48,-9'd66,-9'd53,-9'd46,-9'd61,-9'd74,-9'd101,-9'd98,-9'd73,-9'd41,-9'd5,9'd4,-9'd2,-9'd4,9'd2,9'd3,-9'd1,-9'd2,9'd8,9'd10,9'd16,9'd9,9'd17,9'd47,9'd60,9'd53,9'd22,-9'd20,-9'd54,-9'd59,-9'd42,-9'd18,-9'd15,-9'd25,-9'd42,-9'd64,-9'd60,-9'd38,-9'd6,9'd2,9'd1,9'd0,9'd3,-9'd3,9'd1,-9'd1,-9'd11,-9'd7,-9'd9,9'd7,9'd25,9'd36,9'd24,9'd17,-9'd6,-9'd32,-9'd43,-9'd51,-9'd52,-9'd42,-9'd18,-9'd6,-9'd15,-9'd31,-9'd38,-9'd25,-9'd7,-9'd4,-9'd3,9'd4,-9'd1,-9'd3,9'd4,-9'd6,-9'd25,-9'd38,-9'd33,-9'd10,9'd23,9'd14,9'd6,9'd3,-9'd28,-9'd53,-9'd62,-9'd55,-9'd42,-9'd34,-9'd12,-9'd9,-9'd6,-9'd14,-9'd19,-9'd8,9'd0,-9'd2,-9'd3,9'd4,9'd0,9'd1,-9'd3,-9'd4,-9'd26,-9'd52,-9'd65,-9'd58,-9'd38,-9'd28,-9'd20,-9'd25,-9'd49,-9'd60,-9'd61,-9'd41,-9'd22,-9'd16,9'd0,-9'd5,-9'd7,-9'd1,-9'd6,9'd1,9'd3,-9'd4,-9'd2,-9'd5,9'd3,9'd3,9'd0,-9'd1,-9'd17,-9'd14,-9'd59,-9'd90,-9'd93,-9'd79,-9'd57,-9'd66,-9'd80,-9'd70,-9'd41,-9'd14,9'd0,9'd12,9'd11,9'd1,-9'd1,-9'd5,9'd5,9'd7,-9'd1,9'd1,-9'd4,9'd2,-9'd1,-9'd4,-9'd3,9'd6,9'd12,9'd30,-9'd12,-9'd60,-9'd83,-9'd95,-9'd94,-9'd79,-9'd51,-9'd27,-9'd4,-9'd3,9'd10,9'd9,9'd14,9'd3,9'd10,9'd5,9'd13,9'd9,-9'd1,9'd1,-9'd4,9'd1,9'd2,9'd1,9'd0,9'd6,9'd21,9'd49,9'd22,9'd11,-9'd12,-9'd39,-9'd37,-9'd24,9'd7,9'd8,9'd10,9'd3,9'd7,9'd13,9'd5,9'd2,9'd8,9'd10,9'd18,9'd9,-9'd4,9'd3,-9'd3,-9'd3,-9'd1,-9'd3,-9'd4,-9'd2,9'd19,9'd36,9'd40,9'd50,9'd40,9'd31,9'd28,9'd21,9'd12,-9'd2,9'd0,9'd4,9'd2,9'd11,9'd9,9'd10,9'd7,9'd19,9'd20,9'd1,9'd1,9'd4,9'd4,9'd4,-9'd4,9'd4,9'd0,9'd3,-9'd3,9'd10,9'd21,9'd43,9'd34,9'd27,9'd26,9'd11,-9'd2,-9'd5,9'd5,9'd3,9'd7,9'd4,9'd6,9'd14,9'd26,9'd23,9'd13,9'd0,-9'd4,-9'd1,9'd3,-9'd3,9'd3,-9'd3,-9'd6,9'd3,-9'd1,-9'd6,-9'd8,9'd12,9'd25,9'd17,9'd26,9'd31,9'd26,9'd18,9'd1,9'd13,9'd13,9'd13,9'd15,9'd21,9'd12,9'd12,9'd7,9'd0,9'd2,9'd2,9'd4,-9'd4,9'd1,-9'd3,9'd0,9'd3,-9'd6,-9'd8,-9'd6,9'd10,9'd10,9'd18,9'd29,9'd30,9'd22,9'd17,9'd12,9'd14,9'd4,9'd0,9'd3,9'd6,9'd11,9'd3,-9'd3,9'd2,9'd3,9'd3,9'd1,9'd0,-9'd5,-9'd1,9'd2,-9'd3,-9'd5,-9'd2,-9'd3,-9'd3,9'd4,9'd8,9'd19,9'd24,9'd25,9'd25,9'd17,9'd3,9'd3,9'd6,9'd0,9'd5,9'd6,9'd0,-9'd2,9'd4,9'd4,-9'd2,9'd2,9'd4,-9'd4,-9'd2,9'd4,-9'd1,-9'd1,-9'd2,-9'd1,9'd2,9'd6,9'd0,9'd8,9'd9,9'd11,-9'd1,9'd2,9'd1,9'd1,-9'd5,-9'd2,-9'd3,-9'd1,9'd4,9'd3,9'd2,-9'd4,9'd2,9'd0,-9'd5,-9'd4,9'd1,-9'd1,9'd3,9'd0,-9'd4,-9'd2,9'd0,-9'd2,9'd1,9'd1,9'd0,9'd2,-9'd8,9'd0,-9'd1,-9'd4,-9'd4,9'd0,-9'd1,9'd2,9'd4,9'd1,-9'd1,-9'd3,-9'd3,9'd0,9'd1,-9'd1,-9'd4,-9'd3,9'd3,9'd0,-9'd5,-9'd4,-9'd2,-9'd4,9'd3,9'd4,-9'd1,9'd3,9'd0,-9'd2,-9'd1,-9'd2,-9'd2,9'd3,9'd0,9'd2,9'd2,9'd3,9'd0,9'd0,9'd3,-9'd2};
            // 6
            // weight_bin={9'd0,9'd1,9'd0,-9'd1,9'd2,9'd2,-9'd3,-9'd1,-9'd3,9'd2,9'd1,9'd0,9'd2,9'd0,9'd3,-9'd1,9'd3,9'd2,9'd4,-9'd1,9'd1,-9'd4,9'd4,9'd0,9'd2,-9'd4,-9'd1,9'd4,-9'd2,9'd1,9'd3,9'd2,9'd4,-9'd2,-9'd3,9'd3,9'd1,-9'd2,-9'd2,9'd7,9'd3,9'd8,-9'd2,9'd3,-9'd1,9'd4,9'd5,9'd5,-9'd1,9'd0,-9'd2,-9'd1,9'd1,9'd3,-9'd2,9'd3,-9'd1,9'd0,-9'd3,9'd1,9'd1,9'd3,9'd4,9'd8,9'd9,9'd8,9'd17,9'd19,9'd22,9'd24,9'd20,9'd20,9'd18,9'd22,9'd17,9'd13,9'd11,9'd6,9'd8,9'd6,9'd0,-9'd2,-9'd1,-9'd4,9'd2,9'd3,-9'd3,9'd3,9'd2,-9'd4,9'd5,9'd6,9'd6,9'd13,9'd14,9'd19,9'd22,9'd26,9'd31,9'd31,9'd33,9'd45,9'd46,9'd49,9'd46,9'd43,9'd31,9'd13,9'd8,9'd1,-9'd3,-9'd1,9'd1,-9'd3,9'd0,-9'd4,9'd2,-9'd3,9'd4,9'd4,9'd0,9'd4,9'd2,9'd5,-9'd1,9'd0,9'd2,9'd4,9'd19,9'd37,9'd43,9'd50,9'd47,9'd41,9'd27,9'd20,9'd9,9'd0,-9'd2,9'd3,9'd1,-9'd2,-9'd3,-9'd5,9'd1,-9'd1,-9'd3,-9'd2,-9'd4,9'd1,-9'd2,-9'd24,-9'd24,-9'd30,-9'd25,-9'd22,-9'd9,9'd7,9'd15,9'd33,9'd23,9'd5,-9'd1,-9'd3,9'd0,-9'd3,-9'd2,9'd0,-9'd4,-9'd2,-9'd3,9'd3,-9'd5,-9'd6,-9'd4,-9'd8,-9'd7,-9'd16,-9'd29,-9'd35,-9'd39,-9'd41,-9'd37,-9'd36,-9'd27,-9'd23,-9'd23,-9'd17,-9'd23,-9'd34,-9'd30,-9'd29,-9'd18,-9'd5,-9'd2,9'd2,-9'd1,9'd2,9'd1,9'd3,-9'd7,-9'd10,-9'd10,-9'd13,-9'd19,-9'd23,-9'd30,-9'd32,-9'd45,-9'd51,-9'd46,-9'd36,-9'd42,-9'd47,-9'd60,-9'd69,-9'd66,-9'd60,-9'd56,-9'd38,-9'd15,-9'd10,-9'd1,-9'd1,9'd4,9'd2,-9'd2,-9'd6,-9'd6,-9'd13,-9'd19,-9'd12,-9'd17,-9'd26,-9'd33,-9'd36,-9'd42,-9'd49,-9'd44,-9'd48,-9'd64,-9'd76,-9'd103,-9'd91,-9'd77,-9'd72,-9'd56,-9'd44,-9'd29,-9'd9,-9'd8,-9'd1,-9'd2,-9'd3,-9'd4,-9'd5,-9'd6,-9'd17,-9'd9,-9'd6,9'd1,-9'd13,-9'd23,-9'd21,-9'd21,-9'd31,-9'd31,-9'd53,-9'd83,-9'd98,-9'd104,-9'd80,-9'd68,-9'd59,-9'd52,-9'd38,-9'd24,-9'd14,-9'd6,-9'd2,-9'd3,-9'd3,-9'd2,-9'd4,-9'd5,-9'd6,-9'd4,9'd4,9'd6,-9'd12,-9'd7,-9'd7,-9'd11,-9'd9,-9'd21,-9'd59,-9'd81,-9'd80,-9'd70,-9'd55,-9'd45,-9'd27,-9'd18,-9'd5,-9'd9,-9'd5,9'd2,-9'd4,-9'd3,9'd2,9'd1,9'd1,-9'd2,9'd0,9'd6,9'd11,9'd12,9'd1,9'd3,-9'd4,9'd9,9'd1,-9'd30,-9'd57,-9'd55,-9'd39,-9'd36,-9'd28,-9'd13,9'd7,9'd18,9'd26,9'd6,9'd3,9'd0,9'd0,9'd1,9'd1,-9'd3,-9'd5,-9'd9,9'd0,9'd9,9'd14,9'd2,9'd8,9'd7,9'd12,9'd17,-9'd3,-9'd36,-9'd36,-9'd12,-9'd9,-9'd28,-9'd26,-9'd5,9'd14,9'd35,9'd46,9'd24,-9'd2,-9'd3,9'd3,9'd0,-9'd2,9'd4,9'd2,-9'd4,-9'd1,9'd15,9'd14,9'd4,9'd7,9'd13,9'd21,9'd18,-9'd12,-9'd25,-9'd11,-9'd5,-9'd10,-9'd31,-9'd15,-9'd7,9'd20,9'd47,9'd62,9'd43,9'd6,-9'd5,9'd1,9'd4,9'd2,-9'd4,-9'd5,-9'd11,9'd3,9'd10,9'd9,9'd4,9'd16,9'd29,9'd35,9'd10,-9'd25,-9'd7,9'd13,9'd3,-9'd10,-9'd22,-9'd7,9'd8,9'd30,9'd42,9'd47,9'd29,9'd2,-9'd7,-9'd5,-9'd3,9'd4,9'd4,-9'd7,-9'd17,-9'd5,9'd15,9'd20,9'd8,9'd26,9'd40,9'd48,9'd9,-9'd12,9'd12,9'd18,9'd2,-9'd17,-9'd9,9'd4,9'd12,9'd28,9'd32,9'd28,9'd15,9'd6,-9'd7,-9'd4,-9'd4,9'd3,9'd0,-9'd4,-9'd20,-9'd16,9'd4,9'd23,9'd16,9'd30,9'd58,9'd55,9'd10,-9'd4,9'd12,9'd2,-9'd17,-9'd26,-9'd2,9'd6,9'd7,9'd1,9'd15,9'd16,9'd2,-9'd6,-9'd12,9'd1,9'd3,9'd0,9'd3,-9'd7,-9'd24,-9'd24,-9'd10,9'd15,9'd27,9'd32,9'd62,9'd60,9'd28,9'd9,9'd8,-9'd5,-9'd20,-9'd4,9'd12,9'd12,9'd5,9'd1,9'd2,9'd2,-9'd8,-9'd14,-9'd11,9'd2,9'd1,9'd1,9'd3,-9'd7,-9'd25,-9'd34,-9'd27,9'd2,9'd18,9'd28,9'd52,9'd67,9'd49,9'd17,9'd6,9'd5,9'd16,9'd20,9'd16,9'd17,9'd10,9'd11,9'd4,-9'd10,-9'd20,-9'd11,-9'd7,-9'd3,-9'd4,9'd3,9'd2,-9'd6,-9'd20,-9'd32,-9'd37,-9'd12,9'd11,9'd20,9'd51,9'd67,9'd63,9'd40,9'd21,9'd29,9'd30,9'd22,9'd29,9'd26,9'd8,9'd4,-9'd7,-9'd13,-9'd13,-9'd9,9'd1,-9'd1,9'd0,-9'd3,-9'd3,-9'd5,-9'd19,-9'd28,-9'd35,-9'd33,-9'd15,9'd10,9'd31,9'd40,9'd55,9'd55,9'd53,9'd52,9'd39,9'd28,9'd37,9'd19,9'd8,-9'd14,-9'd16,-9'd12,-9'd11,-9'd1,9'd4,9'd0,9'd1,-9'd1,9'd0,-9'd2,-9'd14,-9'd22,-9'd39,-9'd32,-9'd26,-9'd19,9'd14,9'd31,9'd50,9'd54,9'd62,9'd44,9'd29,9'd22,9'd16,-9'd1,-9'd13,-9'd20,-9'd25,-9'd12,9'd0,9'd3,-9'd1,9'd3,9'd3,9'd3,-9'd2,-9'd2,-9'd7,-9'd16,-9'd22,-9'd37,-9'd46,-9'd35,-9'd30,-9'd26,-9'd17,-9'd4,-9'd15,-9'd4,-9'd8,-9'd20,-9'd30,-9'd27,-9'd28,-9'd23,-9'd12,-9'd10,9'd1,9'd3,9'd3,9'd0,-9'd3,-9'd1,-9'd2,-9'd1,-9'd5,-9'd5,-9'd11,-9'd24,-9'd41,-9'd50,-9'd64,-9'd70,-9'd70,-9'd54,-9'd53,-9'd59,-9'd62,-9'd53,-9'd42,-9'd26,-9'd19,-9'd13,-9'd8,-9'd7,-9'd1,9'd4,9'd4,-9'd3,9'd1,9'd4,9'd0,9'd0,9'd4,-9'd1,-9'd3,-9'd2,-9'd10,-9'd22,-9'd20,-9'd27,-9'd27,-9'd38,-9'd38,-9'd31,-9'd27,-9'd29,-9'd13,-9'd9,-9'd6,-9'd6,-9'd3,9'd2,9'd0,9'd4,-9'd3,-9'd2,-9'd1,9'd2,9'd2,9'd2,-9'd3,-9'd1,9'd1,-9'd4,-9'd1,-9'd3,-9'd4,-9'd5,-9'd5,-9'd13,-9'd11,-9'd6,-9'd10,-9'd6,-9'd6,-9'd3,-9'd3,-9'd3,9'd0,9'd4,9'd0,-9'd1,9'd4,-9'd2,9'd1,9'd0,9'd1,9'd3,9'd1,9'd0,9'd1,9'd0,-9'd2,-9'd1,-9'd4,-9'd1,-9'd5,9'd0,9'd2,-9'd4,-9'd6,9'd2,-9'd4,9'd2,9'd3,-9'd2,9'd0,-9'd2,9'd4,-9'd3,9'd1,-9'd3,9'd4,9'd2,9'd4,-9'd2,9'd2,-9'd4,9'd3,-9'd2,9'd1,9'd2,-9'd3,9'd2,-9'd2,9'd2,-9'd2,9'd0,9'd0,9'd4,9'd1,9'd1,-9'd1,-9'd5,-9'd2,-9'd2,9'd2,9'd0,9'd1,-9'd2};
            // 7
           //  weight_bin={-9'd5,9'd2,9'd2,9'd2,9'd4,-9'd4,9'd1,9'd4,-9'd2,9'd3,9'd2,9'd1,-9'd4,9'd2,9'd4,-9'd1,9'd2,9'd3,-9'd3,-9'd4,9'd2,9'd0,-9'd2,-9'd4,-9'd3,9'd1,-9'd1,-9'd4,9'd0,9'd0,-9'd4,9'd3,9'd5,9'd3,-9'd4,-9'd3,-9'd4,9'd4,-9'd2,9'd3,-9'd2,9'd2,9'd3,-9'd2,9'd2,9'd2,9'd1,-9'd2,-9'd4,9'd1,-9'd4,-9'd2,9'd1,9'd3,9'd3,-9'd4,-9'd2,9'd0,9'd0,-9'd1,-9'd3,-9'd1,-9'd1,-9'd3,9'd1,-9'd4,-9'd4,9'd0,-9'd3,9'd3,-9'd4,-9'd4,9'd3,-9'd1,9'd3,9'd3,9'd4,9'd3,9'd3,-9'd3,-9'd1,9'd0,9'd0,9'd4,9'd1,-9'd4,9'd1,9'd0,9'd2,-9'd2,9'd4,-9'd4,9'd3,9'd3,-9'd6,-9'd7,9'd0,-9'd7,-9'd5,-9'd8,-9'd3,-9'd1,9'd0,9'd1,9'd1,-9'd5,9'd1,9'd4,9'd3,-9'd3,9'd2,9'd1,-9'd3,-9'd4,-9'd3,-9'd4,-9'd2,9'd0,-9'd3,-9'd4,-9'd6,-9'd5,-9'd16,-9'd12,-9'd19,-9'd23,-9'd27,-9'd31,-9'd28,-9'd16,-9'd21,-9'd15,-9'd3,-9'd6,9'd0,-9'd4,-9'd4,-9'd3,9'd0,9'd0,-9'd2,9'd1,9'd3,-9'd2,9'd2,-9'd3,-9'd1,-9'd7,-9'd12,-9'd12,-9'd29,-9'd42,-9'd59,-9'd65,-9'd68,-9'd73,-9'd69,-9'd66,-9'd50,-9'd45,-9'd28,-9'd13,-9'd11,-9'd6,-9'd7,9'd1,-9'd1,9'd3,9'd5,-9'd3,9'd0,-9'd2,9'd3,9'd8,9'd10,9'd17,9'd17,9'd10,9'd3,-9'd12,-9'd34,-9'd59,-9'd60,-9'd50,-9'd36,-9'd35,-9'd31,-9'd34,-9'd35,-9'd18,-9'd22,-9'd12,-9'd8,-9'd2,-9'd4,9'd0,9'd2,9'd3,9'd1,9'd10,9'd13,9'd18,9'd26,9'd40,9'd49,9'd40,9'd32,9'd28,9'd24,9'd1,-9'd3,-9'd6,9'd12,9'd17,9'd14,9'd9,-9'd3,-9'd6,-9'd13,-9'd17,-9'd7,-9'd7,-9'd3,9'd1,9'd1,9'd0,9'd2,9'd10,9'd21,9'd27,9'd31,9'd53,9'd44,9'd30,9'd34,9'd39,9'd37,9'd25,9'd19,9'd23,9'd40,9'd51,9'd41,9'd21,9'd16,-9'd1,-9'd9,-9'd8,-9'd11,-9'd6,-9'd7,-9'd1,9'd0,-9'd2,9'd5,9'd15,9'd27,9'd20,9'd19,9'd29,9'd24,9'd20,9'd29,9'd34,9'd46,9'd38,9'd46,9'd53,9'd67,9'd64,9'd48,9'd41,9'd24,9'd11,9'd0,-9'd12,-9'd12,-9'd9,-9'd3,9'd4,9'd0,9'd1,9'd8,9'd17,9'd21,9'd27,9'd12,9'd7,-9'd1,9'd8,9'd22,9'd24,9'd28,9'd40,9'd53,9'd67,9'd77,9'd70,9'd51,9'd44,9'd34,9'd24,9'd10,-9'd3,-9'd7,-9'd4,-9'd2,-9'd3,-9'd1,9'd2,9'd8,9'd18,9'd26,9'd19,9'd9,9'd4,-9'd4,9'd7,9'd8,9'd4,9'd1,9'd7,9'd3,9'd28,9'd64,9'd54,9'd39,9'd26,9'd23,9'd8,-9'd4,-9'd12,-9'd4,9'd2,-9'd2,9'd3,9'd0,-9'd1,9'd8,9'd18,9'd16,9'd5,-9'd1,9'd0,9'd0,-9'd13,-9'd35,-9'd50,-9'd84,-9'd111,-9'd107,-9'd25,9'd35,9'd29,9'd21,9'd9,-9'd2,-9'd9,-9'd8,-9'd9,-9'd10,9'd2,-9'd4,-9'd2,9'd1,-9'd2,9'd8,9'd13,9'd11,9'd3,-9'd12,-9'd12,-9'd14,-9'd34,-9'd75,-9'd121,-9'd127,-9'd127,-9'd127,-9'd35,9'd13,9'd14,-9'd1,9'd5,-9'd7,-9'd13,-9'd6,-9'd6,-9'd4,9'd1,-9'd2,9'd4,-9'd1,9'd2,9'd7,9'd7,9'd3,-9'd4,-9'd20,-9'd23,-9'd33,-9'd55,-9'd98,-9'd127,-9'd127,-9'd127,-9'd84,-9'd17,9'd10,9'd13,9'd30,9'd23,9'd21,9'd10,9'd12,-9'd4,-9'd6,-9'd3,9'd4,-9'd4,9'd3,9'd4,-9'd2,9'd9,9'd6,-9'd14,-9'd23,-9'd26,-9'd59,-9'd71,-9'd94,-9'd108,-9'd121,-9'd94,-9'd49,-9'd1,9'd7,9'd35,9'd49,9'd44,9'd44,9'd35,9'd15,-9'd4,-9'd6,-9'd3,9'd0,9'd0,9'd1,9'd1,9'd3,9'd3,9'd2,-9'd15,-9'd20,-9'd35,-9'd57,-9'd64,-9'd81,-9'd82,-9'd64,-9'd47,-9'd24,9'd12,9'd15,9'd38,9'd40,9'd41,9'd30,9'd12,-9'd8,-9'd8,-9'd5,9'd0,9'd0,9'd3,9'd4,-9'd3,9'd2,-9'd2,-9'd1,-9'd17,-9'd28,-9'd37,-9'd49,-9'd55,-9'd61,-9'd58,-9'd38,-9'd12,9'd11,9'd7,9'd0,9'd3,9'd12,9'd4,-9'd8,-9'd20,-9'd19,-9'd5,-9'd3,-9'd5,-9'd4,9'd0,9'd3,9'd3,9'd0,9'd0,-9'd13,-9'd22,-9'd40,-9'd50,-9'd54,-9'd55,-9'd66,-9'd50,-9'd20,9'd10,9'd19,9'd0,-9'd13,-9'd14,-9'd17,-9'd27,-9'd32,-9'd34,-9'd27,-9'd15,-9'd8,9'd0,9'd0,9'd3,9'd2,9'd2,9'd3,-9'd2,-9'd14,-9'd30,-9'd49,-9'd49,-9'd58,-9'd63,-9'd53,-9'd43,-9'd18,9'd18,9'd14,-9'd12,-9'd23,-9'd31,-9'd37,-9'd49,-9'd48,-9'd49,-9'd34,-9'd17,-9'd4,-9'd5,-9'd2,9'd3,9'd2,-9'd4,9'd2,9'd0,-9'd14,-9'd28,-9'd47,-9'd57,-9'd62,-9'd56,-9'd41,-9'd29,9'd6,9'd10,9'd9,-9'd18,-9'd34,-9'd49,-9'd55,-9'd56,-9'd57,-9'd47,-9'd36,-9'd18,-9'd8,9'd1,9'd0,-9'd1,9'd2,9'd3,9'd1,-9'd3,-9'd11,-9'd21,-9'd31,-9'd46,-9'd41,-9'd33,-9'd32,-9'd13,-9'd9,9'd1,-9'd3,-9'd18,-9'd30,-9'd43,-9'd58,-9'd53,-9'd46,-9'd36,-9'd30,-9'd14,9'd0,-9'd1,9'd1,-9'd3,9'd1,9'd3,9'd0,-9'd4,-9'd5,-9'd12,-9'd16,-9'd19,-9'd11,-9'd14,-9'd8,-9'd17,-9'd22,-9'd9,-9'd1,-9'd7,-9'd20,-9'd30,-9'd38,-9'd39,-9'd42,-9'd32,-9'd13,-9'd11,9'd0,-9'd5,-9'd1,9'd1,9'd4,-9'd3,-9'd4,-9'd4,9'd2,9'd1,9'd2,9'd13,9'd14,9'd2,9'd8,-9'd1,-9'd10,9'd2,9'd4,9'd11,-9'd5,-9'd5,-9'd18,-9'd28,-9'd25,-9'd16,-9'd11,-9'd10,9'd0,-9'd4,9'd1,-9'd2,-9'd2,9'd0,9'd0,-9'd3,9'd0,9'd18,9'd24,9'd36,9'd36,9'd34,9'd28,9'd21,9'd20,9'd21,9'd20,9'd27,9'd19,9'd15,-9'd5,-9'd11,-9'd18,-9'd10,-9'd12,-9'd10,-9'd4,9'd0,9'd2,-9'd1,-9'd4,9'd0,9'd4,-9'd2,9'd5,9'd14,9'd18,9'd28,9'd42,9'd40,9'd43,9'd50,9'd42,9'd35,9'd42,9'd42,9'd41,9'd33,9'd12,9'd0,-9'd7,-9'd9,-9'd6,-9'd2,-9'd3,9'd2,-9'd1,-9'd1,-9'd4,9'd2,-9'd3,9'd3,9'd0,9'd0,9'd8,9'd10,9'd7,9'd11,9'd14,9'd20,9'd20,9'd21,9'd32,9'd30,9'd28,9'd29,9'd19,9'd8,-9'd4,9'd4,-9'd3,9'd3,9'd4,9'd1,9'd1,-9'd2,9'd1,9'd4,-9'd4,9'd4,-9'd2,9'd1,9'd3,9'd1,-9'd2,-9'd2,9'd2,9'd0,9'd1,9'd2,9'd11,9'd3,9'd5,9'd11,9'd9,9'd7,9'd2,9'd4,-9'd2,9'd2,9'd1,-9'd4,9'd4,9'd2};
            // 8
            // weight_bin={9'd2,9'd3,9'd1,-9'd2,9'd3,9'd0,-9'd2,9'd3,9'd0,9'd1,9'd3,9'd3,9'd0,9'd0,9'd0,9'd2,9'd2,9'd3,-9'd1,-9'd2,-9'd1,9'd3,9'd4,-9'd2,9'd2,9'd4,9'd3,9'd0,-9'd1,9'd4,9'd2,-9'd2,9'd1,-9'd3,-9'd2,9'd4,9'd2,-9'd3,-9'd1,-9'd1,-9'd2,-9'd3,9'd3,9'd3,-9'd2,-9'd5,9'd3,-9'd3,9'd0,-9'd2,-9'd2,9'd3,9'd4,-9'd2,9'd3,-9'd3,-9'd4,9'd1,9'd0,9'd2,9'd3,-9'd2,9'd1,9'd2,9'd0,-9'd1,9'd1,-9'd5,-9'd2,-9'd4,-9'd6,9'd1,-9'd6,-9'd5,9'd1,-9'd5,-9'd2,9'd3,9'd2,9'd2,9'd1,9'd0,9'd4,9'd4,9'd0,-9'd2,-9'd2,9'd0,-9'd4,-9'd4,-9'd5,9'd1,9'd0,-9'd2,-9'd6,-9'd11,-9'd11,-9'd18,-9'd21,-9'd19,-9'd28,-9'd23,-9'd18,-9'd15,-9'd8,-9'd9,9'd0,-9'd1,-9'd3,9'd3,-9'd2,9'd4,-9'd1,9'd4,-9'd3,-9'd1,9'd4,-9'd1,-9'd4,-9'd4,-9'd11,-9'd8,-9'd18,-9'd14,-9'd11,9'd0,9'd3,9'd1,-9'd6,-9'd11,-9'd26,-9'd23,-9'd18,-9'd25,-9'd19,-9'd11,-9'd2,9'd0,9'd4,9'd2,-9'd1,9'd4,-9'd4,-9'd2,-9'd5,9'd0,-9'd6,-9'd11,-9'd21,-9'd12,-9'd22,-9'd3,9'd18,9'd19,9'd25,9'd18,9'd15,9'd15,9'd4,-9'd1,-9'd11,-9'd14,-9'd28,-9'd17,-9'd13,-9'd1,9'd2,9'd0,9'd4,9'd1,-9'd1,-9'd5,-9'd6,-9'd5,-9'd13,-9'd14,-9'd10,-9'd13,-9'd7,-9'd3,9'd6,9'd2,9'd8,9'd22,9'd12,9'd3,9'd1,9'd5,9'd3,9'd3,9'd1,9'd3,9'd1,-9'd3,-9'd3,-9'd4,-9'd2,-9'd1,-9'd4,-9'd5,9'd1,-9'd3,-9'd12,-9'd6,9'd2,-9'd1,-9'd9,-9'd11,-9'd17,-9'd11,-9'd17,-9'd8,-9'd8,-9'd15,9'd1,-9'd10,9'd10,9'd15,9'd9,9'd28,9'd11,-9'd6,-9'd2,-9'd3,-9'd1,9'd1,9'd3,-9'd3,-9'd6,-9'd2,9'd3,9'd11,9'd7,9'd17,9'd0,-9'd3,9'd2,9'd6,-9'd19,-9'd32,-9'd11,-9'd12,9'd1,9'd4,9'd5,9'd14,9'd17,9'd15,9'd11,-9'd13,9'd1,-9'd1,9'd0,9'd0,-9'd1,-9'd2,9'd2,9'd4,9'd15,9'd25,9'd28,9'd22,9'd22,9'd17,9'd11,-9'd9,-9'd44,-9'd55,-9'd38,-9'd22,-9'd6,-9'd2,9'd4,9'd18,9'd30,9'd25,9'd3,-9'd9,9'd0,9'd4,9'd1,9'd4,9'd3,-9'd4,9'd4,9'd10,9'd28,9'd37,9'd38,9'd32,9'd36,9'd17,9'd10,9'd4,-9'd28,-9'd58,-9'd44,-9'd27,-9'd2,9'd8,9'd14,9'd35,9'd45,9'd38,9'd15,9'd8,9'd2,9'd2,9'd3,9'd3,9'd1,-9'd6,9'd7,9'd11,9'd32,9'd43,9'd48,9'd44,9'd26,9'd6,9'd15,9'd38,9'd38,-9'd17,-9'd37,-9'd14,-9'd2,9'd8,9'd31,9'd42,9'd50,9'd41,9'd24,9'd15,9'd3,-9'd1,-9'd4,9'd2,9'd2,9'd2,9'd1,9'd10,9'd13,9'd19,9'd20,9'd24,9'd0,-9'd8,9'd18,9'd56,9'd46,9'd5,-9'd6,-9'd18,-9'd13,9'd6,9'd27,9'd33,9'd29,9'd29,9'd18,9'd4,9'd1,9'd4,-9'd1,9'd3,9'd4,9'd1,-9'd1,-9'd14,-9'd18,-9'd18,-9'd19,-9'd15,-9'd21,-9'd5,9'd35,9'd55,9'd24,9'd21,9'd5,-9'd16,-9'd16,-9'd16,9'd4,9'd1,9'd3,-9'd3,9'd0,-9'd3,-9'd4,-9'd2,9'd1,-9'd4,9'd4,9'd0,-9'd11,-9'd22,-9'd47,-9'd51,-9'd61,-9'd46,-9'd38,9'd9,9'd24,9'd43,9'd27,9'd17,-9'd5,-9'd12,-9'd27,-9'd27,-9'd46,-9'd33,-9'd33,-9'd16,-9'd12,9'd3,9'd3,-9'd4,-9'd2,-9'd2,9'd2,-9'd2,-9'd8,-9'd31,-9'd54,-9'd60,-9'd58,-9'd37,-9'd23,-9'd5,9'd32,9'd38,9'd19,9'd10,-9'd10,-9'd17,-9'd31,-9'd54,-9'd64,-9'd44,-9'd32,-9'd19,-9'd15,-9'd1,-9'd4,9'd3,-9'd1,9'd4,-9'd3,-9'd4,-9'd11,-9'd29,-9'd48,-9'd34,-9'd6,9'd6,9'd4,9'd13,9'd37,9'd25,-9'd3,-9'd4,-9'd12,-9'd29,-9'd41,-9'd52,-9'd48,-9'd48,-9'd35,-9'd14,-9'd12,-9'd4,9'd1,9'd3,9'd3,-9'd2,-9'd5,-9'd2,-9'd14,-9'd28,-9'd34,-9'd5,9'd32,9'd36,9'd21,9'd28,9'd48,9'd19,-9'd15,-9'd22,-9'd17,-9'd34,-9'd39,-9'd30,-9'd23,-9'd29,-9'd24,-9'd10,-9'd12,-9'd9,9'd0,-9'd2,9'd3,9'd2,-9'd2,-9'd10,-9'd24,-9'd26,-9'd19,9'd11,9'd29,9'd45,9'd34,9'd39,9'd32,9'd0,-9'd35,-9'd28,-9'd29,-9'd31,-9'd25,-9'd21,-9'd10,-9'd13,-9'd15,-9'd15,-9'd12,-9'd7,9'd0,9'd1,9'd3,-9'd1,-9'd4,-9'd12,-9'd21,-9'd18,-9'd12,9'd18,9'd27,9'd30,9'd13,9'd1,-9'd1,-9'd33,-9'd45,-9'd26,-9'd20,-9'd22,-9'd12,-9'd11,9'd1,-9'd10,-9'd6,-9'd4,-9'd11,-9'd6,9'd2,9'd4,9'd4,9'd0,-9'd1,-9'd8,-9'd19,-9'd13,-9'd3,9'd19,9'd7,-9'd5,-9'd11,-9'd34,-9'd20,-9'd24,-9'd31,-9'd26,-9'd31,-9'd17,-9'd13,9'd0,-9'd12,9'd3,-9'd3,-9'd3,-9'd14,-9'd5,9'd3,9'd1,-9'd4,-9'd4,-9'd4,-9'd6,-9'd27,-9'd10,-9'd4,9'd16,9'd2,-9'd7,-9'd17,-9'd22,-9'd11,-9'd1,-9'd5,-9'd12,-9'd28,-9'd14,-9'd9,-9'd5,-9'd9,9'd1,9'd0,-9'd11,-9'd11,-9'd4,-9'd5,9'd0,9'd3,-9'd1,9'd2,-9'd7,-9'd21,-9'd27,-9'd12,9'd0,-9'd4,-9'd6,9'd3,9'd17,9'd32,9'd42,9'd29,9'd12,-9'd5,9'd3,9'd10,-9'd6,-9'd8,9'd0,-9'd5,-9'd6,9'd0,-9'd4,9'd1,9'd3,-9'd2,-9'd3,9'd2,-9'd4,-9'd20,-9'd40,-9'd43,-9'd27,-9'd9,-9'd1,9'd10,9'd31,9'd41,9'd59,9'd52,9'd42,9'd35,9'd21,9'd20,9'd19,9'd6,9'd4,-9'd7,9'd0,-9'd3,-9'd4,9'd4,-9'd1,-9'd1,9'd0,9'd3,-9'd3,-9'd10,-9'd23,-9'd35,-9'd37,-9'd18,-9'd14,-9'd3,9'd9,9'd8,9'd13,9'd16,9'd38,9'd31,9'd24,9'd23,9'd27,9'd9,-9'd2,-9'd2,9'd4,-9'd2,9'd1,9'd4,-9'd1,9'd0,9'd1,9'd3,9'd1,-9'd2,-9'd13,-9'd20,-9'd25,-9'd35,-9'd38,-9'd31,-9'd33,-9'd25,-9'd29,-9'd9,-9'd6,-9'd2,-9'd5,-9'd4,9'd2,9'd1,-9'd5,-9'd4,9'd4,9'd2,-9'd5,-9'd1,-9'd1,-9'd2,9'd1,-9'd2,-9'd1,-9'd1,9'd2,-9'd5,-9'd3,-9'd9,-9'd7,-9'd7,-9'd10,-9'd10,-9'd8,-9'd8,-9'd11,-9'd9,-9'd2,-9'd4,-9'd7,-9'd4,9'd1,9'd2,9'd0,9'd3,9'd4,9'd0,9'd3,9'd4,9'd4,9'd5,-9'd3,-9'd2,-9'd2,9'd1,9'd0,9'd0,9'd1,-9'd3,9'd4,-9'd5,9'd2,9'd3,9'd1,9'd3,9'd3,9'd0,9'd2,-9'd1,9'd2,9'd3,9'd3,-9'd3,9'd3,-9'd1,9'd3};
            // 9
            // weight_bin={9'd4,9'd0,-9'd2,-9'd1,9'd2,9'd3,-9'd3,-9'd4,-9'd4,9'd2,9'd3,9'd4,-9'd1,9'd1,9'd1,-9'd1,-9'd3,9'd1,-9'd2,9'd4,9'd3,9'd3,9'd3,9'd0,9'd0,9'd3,-9'd4,9'd2,9'd3,9'd0,9'd1,-9'd4,9'd4,-9'd1,-9'd4,-9'd3,-9'd1,9'd0,-9'd3,-9'd2,9'd3,-9'd2,-9'd4,9'd2,9'd0,9'd1,-9'd3,-9'd4,9'd0,9'd0,-9'd4,-9'd3,9'd1,9'd1,9'd0,9'd1,-9'd4,-9'd1,9'd4,-9'd2,9'd1,9'd1,-9'd3,9'd3,9'd3,9'd4,9'd3,-9'd1,9'd3,9'd0,-9'd5,-9'd4,-9'd5,-9'd3,-9'd6,-9'd3,-9'd5,9'd2,-9'd5,9'd0,-9'd2,9'd0,9'd3,9'd1,-9'd5,-9'd3,-9'd3,9'd1,9'd0,9'd0,9'd3,-9'd3,-9'd3,9'd2,9'd2,9'd1,9'd1,-9'd7,-9'd8,-9'd6,-9'd8,-9'd12,-9'd9,-9'd2,9'd0,-9'd5,-9'd4,9'd3,-9'd4,9'd1,9'd2,9'd0,9'd0,9'd2,9'd2,9'd0,-9'd2,-9'd3,9'd1,9'd1,9'd1,-9'd2,-9'd9,-9'd10,-9'd22,-9'd32,-9'd39,-9'd49,-9'd47,-9'd35,-9'd32,-9'd19,-9'd16,-9'd7,-9'd2,-9'd2,-9'd4,-9'd1,-9'd3,9'd2,9'd2,9'd1,-9'd4,-9'd2,-9'd1,9'd1,-9'd5,-9'd7,-9'd15,-9'd26,-9'd34,-9'd40,-9'd62,-9'd68,-9'd85,-9'd101,-9'd98,-9'd85,-9'd62,-9'd54,-9'd36,-9'd32,-9'd32,-9'd22,-9'd7,-9'd4,9'd2,-9'd2,9'd1,9'd1,-9'd2,-9'd1,-9'd1,-9'd10,-9'd24,-9'd41,-9'd43,-9'd47,-9'd43,-9'd29,-9'd8,9'd9,9'd28,9'd26,9'd10,9'd5,9'd3,-9'd16,-9'd28,-9'd45,-9'd49,-9'd46,-9'd27,-9'd8,9'd1,-9'd3,9'd4,-9'd1,9'd2,9'd0,-9'd16,-9'd25,-9'd43,-9'd52,-9'd52,-9'd42,-9'd21,9'd3,9'd25,9'd45,9'd76,9'd83,9'd64,9'd42,9'd17,-9'd5,-9'd16,-9'd22,-9'd57,-9'd55,-9'd40,-9'd18,9'd0,-9'd4,9'd0,9'd4,9'd2,-9'd6,-9'd23,-9'd39,-9'd41,-9'd53,-9'd31,-9'd24,-9'd18,-9'd9,9'd1,9'd27,9'd51,9'd52,9'd24,9'd2,-9'd3,-9'd15,-9'd21,-9'd19,-9'd41,-9'd48,-9'd33,-9'd19,-9'd7,-9'd3,-9'd4,9'd2,-9'd4,-9'd8,-9'd22,-9'd29,-9'd21,-9'd16,-9'd4,-9'd4,9'd1,9'd7,9'd5,9'd15,9'd30,9'd17,-9'd17,-9'd11,-9'd11,-9'd22,-9'd13,-9'd22,-9'd35,-9'd39,-9'd30,-9'd17,9'd0,-9'd2,-9'd2,-9'd1,-9'd7,-9'd10,-9'd17,-9'd13,9'd7,9'd10,9'd22,9'd15,9'd20,9'd27,9'd11,-9'd15,-9'd13,-9'd31,-9'd26,-9'd1,9'd8,9'd1,9'd13,9'd1,-9'd16,-9'd22,-9'd23,-9'd8,-9'd2,9'd3,9'd0,9'd2,-9'd2,-9'd11,-9'd9,9'd16,9'd37,9'd40,9'd41,9'd24,9'd21,9'd12,-9'd27,-9'd37,-9'd16,-9'd10,9'd1,9'd42,9'd37,9'd41,9'd45,9'd33,9'd10,-9'd6,-9'd9,-9'd3,-9'd3,9'd2,-9'd2,-9'd2,-9'd1,-9'd4,9'd11,9'd33,9'd48,9'd37,9'd33,9'd31,9'd9,-9'd8,-9'd31,9'd11,9'd44,9'd39,9'd30,9'd51,9'd54,9'd65,9'd61,9'd41,9'd11,-9'd6,-9'd13,-9'd5,9'd3,9'd3,9'd0,9'd0,-9'd7,9'd2,9'd12,9'd36,9'd42,9'd23,9'd20,9'd12,9'd3,-9'd21,-9'd10,9'd34,9'd51,9'd39,9'd45,9'd44,9'd58,9'd56,9'd41,9'd18,-9'd12,-9'd25,-9'd19,-9'd7,-9'd3,-9'd2,9'd4,-9'd5,9'd2,9'd4,9'd13,9'd18,9'd23,9'd6,-9'd8,-9'd5,-9'd4,-9'd18,-9'd10,9'd4,9'd2,9'd26,9'd45,9'd50,9'd31,9'd13,-9'd4,-9'd21,-9'd33,-9'd28,-9'd21,-9'd1,9'd2,9'd1,-9'd1,9'd3,-9'd5,-9'd1,9'd7,9'd2,9'd7,9'd1,9'd2,-9'd18,-9'd8,-9'd11,-9'd20,-9'd24,-9'd24,9'd26,9'd45,9'd41,9'd12,-9'd18,-9'd31,-9'd45,-9'd41,-9'd33,-9'd21,-9'd1,-9'd1,-9'd3,9'd4,9'd1,9'd2,-9'd5,-9'd5,9'd0,-9'd9,9'd1,9'd18,9'd3,9'd18,9'd16,-9'd6,-9'd31,-9'd22,9'd15,9'd26,9'd15,-9'd10,-9'd37,-9'd43,-9'd61,-9'd39,-9'd33,-9'd22,-9'd3,-9'd3,9'd4,9'd3,9'd4,9'd0,-9'd9,-9'd8,-9'd20,-9'd23,-9'd2,9'd11,9'd20,9'd24,9'd15,-9'd3,-9'd9,-9'd7,9'd19,9'd2,-9'd7,-9'd27,-9'd42,-9'd41,-9'd48,-9'd36,-9'd28,-9'd17,-9'd3,-9'd3,9'd4,9'd0,-9'd4,9'd0,-9'd10,-9'd16,-9'd32,-9'd41,-9'd32,-9'd19,-9'd2,9'd12,9'd1,-9'd27,-9'd27,-9'd8,9'd8,-9'd11,-9'd18,-9'd31,-9'd20,-9'd31,-9'd35,-9'd27,-9'd27,-9'd17,-9'd3,-9'd2,9'd4,-9'd4,-9'd3,-9'd2,-9'd6,-9'd17,-9'd26,-9'd45,-9'd48,-9'd53,-9'd53,-9'd57,-9'd54,-9'd50,-9'd37,-9'd21,-9'd13,-9'd22,-9'd23,-9'd26,-9'd21,-9'd17,-9'd28,-9'd21,-9'd15,-9'd5,-9'd1,-9'd5,9'd0,9'd3,9'd1,9'd1,-9'd8,-9'd16,-9'd29,-9'd45,-9'd62,-9'd67,-9'd84,-9'd91,-9'd73,-9'd62,-9'd29,-9'd25,-9'd20,-9'd25,-9'd29,-9'd36,-9'd19,-9'd15,-9'd16,-9'd11,-9'd9,9'd2,9'd4,-9'd1,-9'd3,-9'd4,9'd0,-9'd2,9'd1,-9'd10,-9'd21,-9'd37,-9'd52,-9'd67,-9'd68,-9'd72,-9'd64,-9'd42,-9'd35,-9'd24,-9'd33,-9'd35,-9'd45,-9'd39,-9'd21,-9'd9,9'd1,-9'd6,-9'd5,9'd3,-9'd1,-9'd4,-9'd3,-9'd4,9'd0,-9'd4,-9'd1,-9'd10,-9'd16,-9'd28,-9'd46,-9'd42,-9'd41,-9'd38,-9'd42,-9'd32,-9'd41,-9'd42,-9'd50,-9'd44,-9'd44,-9'd39,-9'd14,9'd1,9'd6,9'd4,9'd2,9'd4,9'd3,-9'd4,-9'd3,-9'd1,-9'd2,9'd2,-9'd2,-9'd7,-9'd12,-9'd24,-9'd20,-9'd26,-9'd22,-9'd21,-9'd37,-9'd34,-9'd45,-9'd45,-9'd58,-9'd47,-9'd33,-9'd14,9'd2,9'd19,9'd20,9'd14,9'd12,9'd5,9'd4,-9'd3,-9'd1,9'd3,-9'd3,9'd2,9'd1,-9'd2,-9'd6,-9'd1,9'd3,9'd9,9'd9,9'd3,-9'd12,-9'd13,-9'd27,-9'd30,-9'd29,-9'd10,9'd7,9'd21,9'd31,9'd37,9'd39,9'd24,9'd13,9'd0,-9'd2,-9'd2,9'd3,-9'd1,9'd4,-9'd4,-9'd4,9'd4,9'd8,9'd5,9'd15,9'd32,9'd27,9'd27,9'd23,9'd25,9'd30,9'd22,9'd24,9'd44,9'd57,9'd61,9'd61,9'd51,9'd38,9'd16,9'd7,9'd4,-9'd3,9'd4,9'd0,-9'd4,9'd2,9'd2,-9'd1,9'd0,-9'd1,9'd11,9'd10,9'd12,9'd20,9'd22,9'd23,9'd26,9'd32,9'd38,9'd20,9'd18,9'd16,9'd22,9'd18,9'd14,9'd11,9'd5,9'd3,-9'd2,-9'd2,-9'd3,9'd1,-9'd3,9'd1,9'd0,-9'd1,-9'd1,-9'd3,-9'd4,9'd3,-9'd2,-9'd1,-9'd3,9'd0,-9'd4,-9'd1,-9'd3,9'd0,9'd2,-9'd7,9'd1,-9'd3,9'd3,-9'd4,9'd3,9'd2,9'd4,9'd1,9'd0,-9'd3};
            ///

            #5;
	    @(negedge clk);
                rst_n = 1;
	       
	    #5;
	    @(negedge clk);
	    	enable = 1;
	    
	    // Logic for program termination
            @(negedge finish)
	        $display("Finishing the run!");
            
	    #20;

            //prajyotg: Writing data into file
            $fdisplay(write_data, "%0d",product);

            $fclose("write_out.txt");

            $finish;
    end
endmodule

//prajyotg :: extra input samples
//        if(product != {13'd30,13'd36,13'd42,13'd66,13'd81,13'd96,13'd90,13'd111,13'd132}) begin   
//            $display("test 1 SUCCESS");
//        end else begin
//            $display("test 2 FAILED");
//        end

	    //input_bin = {4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4};
	    //weight_bin = {4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1, 4'd1};
        //#30;
        //if(product == {13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12, 13'd12}) begin 
        //    $display("test 2 SUCCESS");
        //end else begin
        //    $display("test 2 FAILED");
        //end
	    //@(posedge clk);
            // for (i=0; i<50; i=i+1)
   	    // 	@(posedge clk) ; 
